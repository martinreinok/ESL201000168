// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H7YP(K8PDO?D?0)4<EV4-R9MRC<'DGB'%M.FF5G9]"7BB;3W4W"!4SP  
H\[P$/NK1Y6D87=V043"!N@4(XON*X:H_Q@_O8L#FZJZ]4XK6/4EXC   
HPL\ +&HM67(6>.?2/_%WT,#GR_1I9?4A\3R,^M"/7WJZ4MC^(4I@-@  
H[D0L[W!,ZG2/2?JG6FO$"7)M32 =BP\7^&BHEH)/^@MI W/J ;TTR0  
HXXKUKO=4//Z.F)^6N W?'@,H.O4_S4[OS'4=JXFZIY; CZP-781R:P  
`pragma protect encoding=(enctype="uuencode",bytes=17984       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@7QNM29\)QV8$)/M3PKIS[GC?U-WQQGVT;5\+BUGS[&L 
@\496<OQB>B\CO ZLE!*1+>CH0;H/-C[!Y#!NJ:Q5P?  
@;P!V,\3>L;NK[M% B#]1D%08\X+53]'W9$D*V^>GT>H 
@%F2-)*'Q@_<N:^D=])"QZ=LQVZ'/_G\4_G:IR]M0!7L 
@<3 =B3CF395/7-@=U>%15F \8C?VEG#4ILO)N]*:%E0 
@8:&%R%GER.I9!+GCD!V'$:PO2;@X<9:G*2=29E+;M84 
@\B"&CX"6<_%/8*_>P1:79CV;%0_=DK3(W,;X:'\:Z'T 
@'IX#I3RX#L27,5A;'N9K()84<K.?588N=4'IRS ^Y+P 
@D((@$@35K&E>,N.!];R5FF7-[+V0FIIH7XZKA+RV[H8 
@93,6;!]1MU+THIB2 UQ>MHE]\R3CL=W&<$UH"A<5E4  
@=& ^]335/[9"A/'&/B H"C!F9+_AU15W*XMT0%(W=[\ 
@CL()OQ KN!*Z )C3Y][MH5#.[P775[I\XPZ="66?Q78 
@IX\+-E:U63@MZSWJ?9 >.EW?I 2.H!-TPAF)&-KL \4 
@&0?3CJ6J9,U@ UB$!8']K"AW@_ 1-;H7X/#<E+)D=;, 
@!ZT3*S:-[=1 '84X".DQS"RA45^!%1>BY]H(;CY[_'@ 
@31K2:1?@K=58@$)-#BOK(1QD'2'.O&.T-)-R(@=3)(( 
@]-;C1T6JY/G$6:\%<C,).B/=@ZT*OU-29_= F32S7V\ 
@S&6!KB<TFR+VGD>*@\RM,_HP=MN$ U]6&]X%):3A''L 
@+Z:JG$F=65@.ZSQSO#_#4"BHQ(A/F34W)BO1'D<=B%$ 
@=?-Y[S==<%/YIE=SK%I[K'!@4OV%$A^7V+:C>Y6:IL$ 
@)!)_EP4,J4W#, 1< )_;Q'XR<E>G%1N$I"H>(BX^RU8 
@%(<R)?R3AWY$'LG7XUUK;SJKX5G@<F:6_I>B:W[$*$, 
@.'%]O$9"FL.&M? =PN?FRRU,C,]X_(;*ZJ,QBC>YC&< 
@O#!IY($1A /U=;(!@1"]P6%D+XXX/!)>O$5!@IVR89$ 
@*>"K4ZJ\K-&G]P'UD50@^*ENZ@M81-IF9K4+G=_;K., 
@CM)D&6$6*L!_B8R4?]Y4Z,#%!9Y@O%>*W,4N+EQ=!5  
@Z>3SRLO(_8\N@OM-PTWNUV9V:?F.I:KX;9KZG_)&LM( 
@HD/,Q$6[\\B[=9$$$>'FJ5QM2^I)6[51%GN3USD'1?T 
@6Z#6_N\=1G<<C8)5W%YF:Q42(6P\W?)9\6PF<E2_L!8 
@ OO/6$%IGS <^<9&M.ZGQR/!^%+C9<;!-O#UXFM;UI< 
@1X_*2#XWC/1X[1I9.T4-3I$CY&U:IF; W+>>![ .<;@ 
@(>TG;AG1*'-Y%"*L/2H^TT8V49>6V%TW*<T$4E5B#,  
@5;Y*_?U[!N%I_\3M]T!3,/5%,*R_GN8RD'-44=FE>&, 
@LNM*?].4I9^]538-/&K590G=2;)H4/2&K,"K56JD)F8 
@!_S8*@'KE#G,*T=T'Z\G-]JP+EO#J0\CY 6-G?7UI < 
@\;M!5!_:&2@*T'PW]IA"UDYI9QPYA/KO[00?AV @O>( 
@F5-349C!!;3K85J0% 7%0-\>V9%46G1[>?E9K5(B/?P 
@+.TGHF34K",Y! Z\Y@70BHAT)%/%<D/&#<UB'Z(WUYL 
@B^ S!W7,4;V('LY(@Y#@;8B/C=D.)()'T;'#:7<BGF@ 
@%R-*4ES2FE<=CTN;B>+W69L/,VR%I_2$*_.;0BLAJ^, 
@BAA6T()RGKD(&))4(M]N?NL]M*WX,PLG<:DE7\HT0)D 
@:-F-DD9%6T-F*[_; TZGS4$_<;\9_V@FUH<D@H<?5>0 
@X.J4C[ZO($)G2J&TL/O]:;W3H_2^5?$DT)>S_4U+?90 
@X?,S'/2M*]%A3)B#^4++(\DT*6&:N[]^O_E>W17U50$ 
@#("+#*_$W_K:KQK=* AG4ZP>;9A&PX?>_GVKWC=H ]8 
@1S+7I>?J-R(=4.5,NXQZ$#7&S]!YR;;:%!BR4:XN4>0 
@O(U\D.]UY;I_7K?XC_8EN;<U8S]6,[7.^CBQ)UO-Z04 
@5@]E8>I+'"S!X],QPKYCE.>"T"A7'1)^O??<L!$GI9D 
@X8?NZRNEDA*R<!=L_T A\7X8GG8M\$[*+OU 35(>:B4 
@<F[#G4=63"P$9;R=^ *'R:*D!7&=4VE>FSD)S!2[$"H 
@'L-<& AZ#,S#A<LU!4RSO2V5>D\<IT5-.PMFI75@)V( 
@<&%12%5#$6W^L7,\JS6\)+ 30]Z9T,VVWZ+S K\1IN4 
@/1.6? J#U"O UG+I00Y7]D<;:;?4L>T).;[P;G37L=H 
@'RE0.H38=*%R$8-E6N6*/#1V835M].%6S;I^NXRTT4D 
@E;35D@W>.6"HS:PXN=3 +=Y+GK_<PSL']].'J4QF.*L 
@3?C,("1/&=L'/O^=+NYCK-CZ/.2$$]^CW"MXGCAN_:4 
@^SPOZY_-8(UBO2N8-/^EUKD(>/)Y4$)I8O#6N'0 @M, 
@]C.E6F5DI2"%@$5@.\D2@FK *^K:K&-=9LT+5US0G]0 
@LSZ8_M/Z,8RKH ?9$(V2$XF><MU3*+Q3I9\]J'!PT,L 
@>)!C2<N-EK6JS%%QO6WL33@X\Q/N2:5( YG"P16 R>H 
@[-0X>[9^HQ)3O)I69?!P+VJ4KK7#Y+J<HOCRI,F;RB< 
@'_PO]Z.SP01B[JQT5PL5@VJ[KR_B/RF/'!($N*24;B\ 
@5]&5"%M9Z)RA)6PG9A/;]M=+&6!&#$=I"'3L+*P ;-( 
@J5<=8^W=:[)OP98T[HO&9&\FO03;'O;SY><:KP1J;8\ 
@'D9DD A:XQXN.@J&A,8*>/O[]1I+GRJE#S]7DU+OH^T 
@?]+4<2O50?B'][?NUC"DFCBKM%)X5-Q_+1,JB"NMHW< 
@O5,3.4? ,09Z<<X6C"QHE*,9?7I.3GGWZXNA&8,7+ T 
@MI:<ZQ@+X[3#G@;,%\<GW.>K%A? R6+**5OHFB+]D&X 
@OV8=KW5]_P]0A(M4;TT7E^1D3W1U,V)E<XO->M"D%Q4 
@6WD.MZC^%K&SS2?@UFU[.3PM)&\'EI=5A5)(4">?UGT 
@]1".M[M"8-U2P?M"<>@-?/07-=C[3M?>#_8SA/&!( L 
@"P$_Y0O*040]M*[0P+0^O9M5@K=!Q)<_9#]LU=ZF,P0 
@8)B'I%W-)3+=;4/Q\O0WT#]L'(E )9ELZ$U);[ VDXP 
@ \(9=[7CDDC4714??<M8H>!$%AK)FS*@_!%3$V?0,6L 
@(%-%T&[V90F-8>1O']^L5HJ&>$(XO>'.5])?YX?=<TL 
@(-<;)^X\<1S>*,1SQ5%:(,(?\636"KISA;%P7QK<<L4 
@0UIILB]Y,MQ9;*B5(M>FZOM@GJ0\_B$$%OJ"SYP#+9  
@1*LM[<4T= O:+>2:246-QM^3AVZBVQT9(IU3)[#WT/\ 
@V^C_7D3:U<Y=-$'P3580YH7FD62SU8GCB(]NF[ZS*<D 
@!<#,&9RN+:*E48G:MZE ?*J<O>U8D2%'\L,NQ0(^#C@ 
@Y\]PW&N>.X!6Y=MSF)OG2]U29IIEH@#*37KP]9X6)6$ 
@#K^SPY6@KZQ9KRM1#9@$Z$)4?F[9M"YL%)*II\,QXAD 
@A:)4(KYJ6R;7UN*0UY)#U&IH1M>Z*;K".&M#&N7Y")H 
@'Y8D[A,%)@R*I<B5(-!9Z7!LAJR/AZF<PG>@Z/'6+7  
@QJ]]$[,(.C''BCX7IPE'.*,\VX#[<U"GME*'],)%FLL 
@K>]!1J>XX4*#]C1T,K>][B+P72R(QCHLTU]$<SIAD9T 
@8%.PM!A+V,,2@R0H=Y(JF0UDXMJ.'&/++.A!'ZK5_"  
@P##EC0C_Y9X,G'$R:V#EJ-#ZVF,E<I++/_LILCR'L*< 
@ Y['G])%;2@D</64T8?I+570R7QB6?6^H[K%$0!#;ZT 
@G*G DO<7*_AOEE/[8[-EQ XV5/YO_D"P>ZGEV_+RAMH 
@CN\4S&WX 123G2M!MY9=V6WY8+UO[-7#7[Z-ZNO>-Q< 
@2 QM)CAR\%]6 9KGFKJZ@7M(V0''*@9<M'%$'_%X-5X 
@TXN0@--G>?#[01N.?X.H&V!E]RM$M!N]EB VI+LL&D  
@*GXELE-33P"+*=32+LQ;  -1U2\3HO:LK< XN4X9>,8 
@GR]^:#,F&:>*U].O5T<9EU9'.1\CZ>1D;OQ3A+GXS-@ 
@VJ%)+ACV.=A34U>%D9I4+!=(C/Y!/R-=H\.)>2NR0$8 
@B<"'P&.8[(D73T2BN$+6]0=/V8LWS6']"#/&$;WON<8 
@;7NOBG<7$20)^YQO;Q>VV&0HH@Z_SOT_#;H(I1N<>]\ 
@FM.T!Q*BO\%J8%Z(8_-0Q0+?%:RT1=C0KT\^*48,O;\ 
@2(B*U;M<.;\ 957CFIF\J/S^[W1NB&70>O1U(-MIAV8 
@G-@?\A-F?\:'2QOSDOK=LX_R%=-B3*1X@$DM9-.'BMD 
@/Q\O9Y<.5HHEJHMA2O22I+$E7C,+JFS@D 1/ 3LO.<P 
@A<DM*F:CO&IS+7ZP2HWHQ#+A^^.0IZ+FF@R\+* 0L-\ 
@3AAD:Y%(4 Z" T2RRB=0\,%"3;=@A= 3B:$:@SSA>^\ 
@NJFP\W(9Y:7U+:Z]TW)N\DT=" U8#76GX?Y4Y4RF^K4 
@=%G+A+1-]@++$QI7 'F#UY07K1W$F&TNV&H[SN\^V_$ 
@ 2Z_9 ZQ6C*$X799+1B ]JW,-0#[DE1'(K8[),$+L-8 
@UPWBSWC7_H R-Z\?M6$55N].%W>/4F604"J'X%?7ALT 
@D?R..R/=PNE>9_&[T'C1U3RXL(KU-7CUH<D[%/P@*"L 
@,XM><G4M%:..J>-CW^T3G^8$4WOL9[HGDJ,&M5+XJ<< 
@)T),D:++^'*L945P!!;_ S>@,#B!@,XL\@J:P]+T@:$ 
@!=Y0]Y(3L3>6.&FX@\7R4*1JAYC#ATLC%XPR6:,Z)I  
@#\J)7G,K 5@E*"<4VC%9<'OGB $] LIII7"]7 5W]1$ 
@\<9SU:$P@?$]425'T,I>Y5[9)EA$U6E?&>1^;3B,:J$ 
@^"@M_:H33V6T(#C.3@N-4!-;\Y1&]4?H03VQ!O$)D14 
@=S^,4["Q\V? 6F#W2K[/3D0J"1B"QF!Q>/ $'.Q1" < 
@>1X?93)L#J9:,RH:% :&.4/GR;EA/3?ZF7FF03.&)>( 
@X]SA(>/8K+UU[Z=$A@]U(1TNX,U%VC[,B3-.#S\D#%P 
@UJBV3L=QOZ\Y8<AQ+U_8=F[D86DC-J7KL91KR-6&^,  
@ 0LAIOP^-@"4H"#LM?^N#>4L$)#5(-(B5WAJ6C=&CHH 
@9 1*H3* #!B+KE6#@9"ZC736/AP*B5C.6I$[!,MOME, 
@W)".<^JP.,X5*1  KRB&@H6V6Q*'$FE963/V2HJFD8\ 
@]6'3>/+53$B W0S.D_32DLJJ?ZN >OZ\8@UTNMN:74\ 
@8>IST-523KU_$R2+DAOG =N.L->1$<_Z2Z&XCSS7WBH 
@;XQ<,Y<%V@3$#C\V<]/[.)5!A+0Y(57*:!\@@9"Y"Z8 
@9S$$. :.Q7;*#M9U.E:V_8V_R.6! #]1*>&6LPE:_6, 
@7B*-"F;CDGZEW'?S"]>Q@CS4./QUY>8_R_/[.1QI/P\ 
@)FS]Z/OTU3409?/%M^[K^1O.:S'3NQ<[HUD"3X?\7S@ 
@_DST.KHD(0^B;+X9R H6A8;G<9U!MT"#+J ;22/X@<4 
@N:7#E/O:MQ"TPNM5>[!JVJ)VQVX5;;M2[5H1$?S!<H( 
@N/OGUR H#_T;)R><1=FYKU"?]B>$P1[;1DSZ!PTQF=X 
@'YWO%H%"R[#&_-DYYT0L.16>%G9V)H\ ?LO,!W*WH#T 
@P:0@''=C6=K?IR*\Z3Q%DPRBF&Z58]% B&8M \_W[%$ 
@G8_/\8BS#N$H]E"O229,(+?^I@$!!#&".K;6 Q!=F=@ 
@>R/V 31!BU/4-Z&<4I4K2E/A'P.L;JY%6#;I_J1(E%  
@AV;V7VF#]T@T<P;=I9A!B<G=M_!+ V^D*4BP2[Y?ISP 
@_A_T\@?,#JL/%+"ATF[I=;KQAJXC!7WUL6FYVP)K0%8 
@8SB3/&OY/B6JV#NO?*;!Y5C2%_MBBY4-D:,;OZ&YZUL 
@*;ON46"S^@*E^1PNZ80CY^LUY;ACL2+2HLC\^:: D>8 
@=Q:B:XRR;;UJ=-@NLE/.TRPQI+4D':D'9X:^J&(BP1< 
@-(JKO0M(_?6>4"\E"0ICCR'H8SWBG0=0B7NE!M<CYB8 
@B.A$QV$V#_&J#V K9-.2SND,_8N?SSV_Q3.F*][F=G  
@5=Q)'\,F55YR<2T0/5CG*"CSSO5)_3?Y.DDV+['&$G( 
@S*!?J)<E6]2<$@AWZ)'JP[[88W@M*V#LO:L7YP^-1'L 
@'>Q0+VGPAM(?.I4VF'%')T]FYR&5KZ3ILV.O]T$-LVH 
@=QL1<MG"'+"]O3'2&*PZD4/+U+0UP7DN"R"A->[EJ=8 
@K 7_/-T#Z^,.&/5]6DK:]\BX+D+D%K'6JSSP+I<:D90 
@D]&4V:$0LV)BQ#Q <"7@1 WI"44<$"PQKB.!N"7Z\U< 
@#KE-R*=8"#6A(Y;T& V>5A2 "/Q=-,;G?OZJ0XKM*+$ 
@R]S(#!.2?E^/83SW.1YB)UK2@4HF9,W@6U[6Y$)N3;< 
@+=WEXSK?7. ^#N$4*H7N!8;2M7,N8552F7(V#84 */$ 
@4$G^?YL1"P-*LM?).W?0\)#G;M:BWF:0>\J-1B!RH6D 
@FY>CMU,)5/:S+O/AS^KL@@&-$Q7)?D%@=HV,3QJ^8.D 
@7'B2F)_HS#)9(+:P:E&Y,SSIH!0 "\!8V+)1*8,0TZ< 
@JA5[2&L4W2:Y4Q)_,J;-CR5@Y?@_?,K]$AY90"S_\I@ 
@P=^]^24[AIML--X I?G/2?AG_GZ'K)%W$C2ITW(0#($ 
@Z2[0NAR8SY=38-8]S;XA9+2X+G&26M3?PL,K-42"HY8 
@O;)+2GDQAWM!FJS PR^ER.+\ZRM>45[#*ZO[6;];N.@ 
@36 -_U01QF#2?9EHJB( DW_=!G+',<AC :\7V:^6W:D 
@U%I#C22I;7:=@_I@C]/?.G5@8ER7P0"D* "7Z'K:ETP 
@(V'SM2H@)O2<9075NGS+F%\^RH]2JN*?_O]!,[ UYLH 
@J.\?:@CP02MM ?+;:.3B' \$AM^;898QL8>JI)T6 X\ 
@U%4XNV!AI?KS[(NF6VH_R!B.^UH@8X%YNXX(F;MR&[  
@GJ/M/(??'/1</DVZ('E.7S(J7L &9?&/111O!["KU;\ 
@,S:W^"7==0]7L0UB^?D)2*SJ:4"(H-+<Y*)0'_+PV!X 
@1X/P&^D ,@>?ORZ=RSRJ^UI%#'G]9J_3'<_\@3TEFRP 
@6$- A3B7I-#%'JTP.[BS&LFCO,0"W"-QY%K;9JJ1,QH 
@!"H/49_DW'$/17C]/%5PB5]6J1U6230]]Q=W=.W)1MH 
@:?S)*#BR;H/(;JW'X>R,LZ$*,G7I%S4T8V2^>[ BV<X 
@LK"U2^(N!>+EFBF"<53):%=WW,&+)J(B3I4 XI>XNC\ 
@O&@#/8RRZA 6GVA71#7%5[XU:\V$1)+463SLJ2ND^\0 
@I<1[?DK5"?;=(([#F, \8\8/!P:(+#=4ID2.O54'C"0 
@,1IY6F5"NX/E[S')QX(Q8%]?<Y^]C;9L!Z\\0*<IZ.\ 
@980!19]I0+BP'V%QVFY#S&N$HB/AY+7JG9ZQ:OUORZ@ 
@IATV\L^<A:R^@#5P>L&IVU<_.@J)+R_O.QJ$,1<1'^< 
@Z#;L>#ZRO*JGKPFH,@*$5<JI-K[H,VTH?0Q0;GC%"\0 
@1:45B!#?-%?<%+@#M(09\D?S1-7XMZD<<QC-**'46W, 
@4TZH;R$XB<ZO >R_']:RN6*1%['GEP>LJ66-0]&:3KT 
@]<S%[G%0-7$4W>7%:\PXJSC)L&=\M_\=\'D>^0=@2EL 
@SPA'&L)F/68Q(=,Q&0!!^(BNK:L=Z<(T"OEQOFS%@4$ 
@4V/%$K\=TJ#S%^A%PLH*U"=B8<YV8[O9RN.4(FL+#1T 
@ <@PB_"YHWL@GWOH9RFG$#X)-Y5X/1,XK<.MA93$%W\ 
@-_Q78#,<Q[O\X-9# 8=F"%!K*P>7IBX+J<?_4.SJ(60 
@TYF-]%C16:@8B/B*JE:0PSI?MJ,WI N1PA8.ONU@+ML 
@)<<4N))0HD6.#SM/H"4_>0.@#U&Q3A?EM.'C??,QZ$X 
@TN/8N\T3USQ,!ZNYHZ_0N"&%U3<H/MZA'<*R1 KOT+< 
@^;W76:+PTVKH\[%B((+JH6>+G(U;;,B  K2:G9S"AG  
@"^0-JO%-@+]FP8XX]G64"H#DPZZTE$JU1Q!PM/!-ED, 
@+OIH"/E;$@RG5HC*B!"(,'01(HZ('E>#$*"CXR0<"&@ 
@<[/?YKB].[TTZ%XK(QDB6/[51,R1LJ>([+.F<?<'XBT 
@S9MZGV-1YHF=&STE>W.<M$CU!,SA5J)AG&+1?*E7EF  
@1DCP8]$0R2?5P)>D9[80.5=[DN Q[_/U1D&(YE]:@=  
@Z)WX7V$;H8ZF#$:S(+$1EEFD1!QA=CY)@$Y'_M#5&R@ 
@R/]-R4;5DS7/Y>(&E_(/RRRH7WHDT( SKDE(\#@Z4ZL 
@'9@2?8%,T;NGUK4DOFF*2&P8(ZH:+8_/EHJH3?4.+#P 
@?)O1I"GB@JQJW73Y4IQX)D'03(ZE88Y@Y-16:;2"9E  
@^0H>C+.N$7P1'R/-5#Q"J\+ESD,GTEX:5"2F.L%(T&H 
@PRZ#[JXI!/'[;D^[Q210;UM/VEA Z^2POCJK>?OJQ34 
@Z_J40W3&L?;]5D^&14-W/6AY?-=W7$SY.?@H?2-(X)< 
@5K1#B -7OY\K.!-VH4GD='36W\>.2RV;7?I@UP'%2N0 
@6>@/>7^6L!P>WQ(&WQJ@8RAEY^TPHC:,S4%^(E70,ZX 
@13J4UEU/NB9%#%,S$=V<_TEV%RY)B4OXT:2Q2.OL9V  
@23@6Q.:XHKHV5*F66W2QA'KEJZG]>2G2MQWI_Y!5VU0 
@!9/Y58/TE7 +TW8Y+6&).#$)(/Q[*4#5^=?;_B?1>+, 
@+9BG;$&Z4F _>@,@"2B1BK'.MQ3<Y@N)N>4ORG>3.DH 
@6.AE=+ZH>Q Y>NX]SZ*ADKF^\Z#4A\#ZA+GL+E[D4AL 
@B]')_@@X1PRJ2WB0=A'F#U?1 ;1 $#J$,'!'$]*PB7, 
@3%-O>B=5UYC2&UGDHT,NOYP3K+GLG8^1BWGH9QB)>;4 
@M-4*LQIY2#<G8!,6[SC]%B.EO:#3);'&F0-#\MC&_Y@ 
@Y1E2Z\7KOOVAOC6YN<YR+>C$Q6QZL^8[!?R,H]53G4P 
@+VON$3CF49]*!\,Y@QOV0CR*"52)MB]-'"GP>A&@3*D 
@C/,8GF3,#&9(5[K(;M5F._,=P!1C4XFYF<B-L]15:,T 
@T>UT;9I!=V6V'8)1I-JG\QF&Q!C\3N9ZX[EAR4J 4KT 
@25X>1!JZM$/9FU> ]+](YLB)Y\/-ZC;MY#T08/S04@T 
@]^02T.]52Y#8E6/&#-4?"[:C7P2Y1ZI)R005MT7^W\4 
@)T798LG/Q@M_R]PI&.L(>_=M<G;JW1YG NK5(C#NN@< 
@)DXR]0'O(W3G #N).=-J@*RYB^93<1Z(Z_?+6>+9F_\ 
@M/<$V_O]3-B^*=0".FAU#DGW.EM'Y##FC)7NQ8,I.?< 
@ST%P,5OH*GR&\E["%ZS>2)8><:.>N>TA>M=H;HN #?0 
@'A/@VH6'1JWC<-WK)GK=?YT\*!!=2= 0#<T,=1Q0!XP 
@8(6.]&NQ^"?G@2O?(7]A=.,=!0'N/:-G<S <J,06^_( 
@1+& 8:GGP&[XF%.#7EF4'LM91Z6LF3,M'((P5KM* $X 
@@"1.- O1/JJX.]$:T.(X>DMIWQI_@OY?'C]5@CM5OYD 
@J'V$VA5RU1WJPN>_]AW9RZ?^DB-*RH."DY5L/="0G5, 
@X?"*8UK_)<&B9[88#P#=:$T>?P,B)6U=Z"D<K?&NW), 
@J\:T2W?^,?#%??+W14!;%<8$Y_]2>^&!AYJ4O)+'@NT 
@F!2Q.(!2W@,Q'O,E;P)'GE1F?1P-8:S-W#'1LGM-H_8 
@@ >$$U]I%UYT?)W<R%8@M[/LT5]];#CLDI8U+B. 2Z4 
@KJN$9+/GG+PJ3>@E0E734BAZ"#G=O=7/V_-J![-]&3( 
@!9+QE*9W'#H.Z>\WK'UHG;D%/]3,\T<LW[+R?&&CZL( 
@0@2Z:''Y@,8Y5+&_I"8!!E3W0C@GPY)3GTQE8_'B2;0 
@Y#4'#V"M"K6!\_W6M83XY+HN)EHK&1Q@"!R>( [0M-X 
@^/]R&AZIH]6.G5V=1W08P56GUD\>>'=ND\=%Z%Y(W?H 
@\DIB. G&MX^\>2$77@>.!M1+;ZRB?JGZ76^U:F]'.?X 
@)E\J*&C5=YK]_S7(74BRSWV;SNE&"]56'T=N ;/:S)@ 
@=:-,F-*](P4RO:6[N>F\K5_'Z(--;5YH@'4Z'#/3;FP 
@?5 Z1)8$WYWQ<[<;Z 'M+G:"<*ID"E:"2F%K U/4=., 
@]KB_$+FJ'RTI ZDSC77GC+K?P*)WCSS6_1R/5&J.5(  
@5I-YBF>-6A)U:\?SVN8^$ \?&KL,H=U6R5^JI7&PR&( 
@26JCZ.BXC' B=W\H[MU,)5 >N,QX@R:]<&*%X7>=:O( 
@Q%(9H*.RJ3?B*T7_RJ+92:-Q2P)JM.XA=LOR9DD8>.  
@)_U]V:G%&ER=QH+Q5;A_24T^4"HUV XM:5Z1T3]]/*$ 
@YMB1K\W3%]7@8$TZ@R,@+7744CO</;<L-KW.Y5P45&0 
@-WQ-*O?VK5*7ODV,S'R-\;"'CF5]T+?:\Z\74FO(/6$ 
@850]]9*L=BY6W(KA>VOD*<Z4+A\G;6*'!1UX+HS-T8  
@8EXUM8Z(^X(C[!G2F=B,#@*48TP BF7O5\CN;?.)!+D 
@=\XM0FA(GE_1@GD1O=0E4[;E/;(F>T)'D407^KNBG2@ 
@&IRSH\T:M6?9>%&RXH.#=%8Z-5O+^88H"MO:"8C%T$P 
@ERAM-M#,AKT'X=SS^*8ZXRL?"&D[J%@W#P0V6\BD<HD 
@^[+-.P%@%,?:YH7$?$6C>DWP:T<D*GBQ@F3N U+-O64 
@\LR@HR/GKN('[F_1 Z\Z"7>,F#&MYF(?\/ORBPCCVJ4 
@4Z]&7'B)#W_F\(M:9^K!^#O\[,0OF^P_6=+,EIN>]1, 
@<2,]E0'F.4?@%H(#<M=:GZX;C'3D/T?()AJ%^H&?K\T 
@%0!3N43,W?#[42E<)*]+[]%9QX=+6?^3U(<PW<:G.5\ 
@,=%? ]=/#Y)>2(\S@DWP-:__W.GX.\::'9HW[![=,^< 
@C]PYFX!'=HU+^5P,4A;VP:\_^*TTGAM3\GC/N8,)G,$ 
@A*&(5*B!G @N<TV:3G08#YTA9RSQUX*8GV">T8W%I9L 
@#<<*OQ]MXH'3)K" XU1VT@$[A?Q74;O]\2;J>?&;[90 
@V.JB\)7")8A<2P>E_%+M7-J^O4I]VI>!<CXTV]G0*$H 
@12MY_5.R(DZD\(^^9EVKD9SH8YJ^LC^@V,IF<U)+R]L 
@;=NSJ^4X)B^$EZFH,3J\M&[0% F83MP;L1&#HGU@2I8 
@(]O;(]<U[[JL0ED!>8K7.C]R8%]_);FKC * [_E#A', 
@4F%T<=> 4%/KH5-&S[&^YKC!4W^XTG=A#OV_F(K\]O< 
@ ?._2L$89(B=98QC*4*)^$X#\;8F9XJC;.*TN9DBGJ0 
@I+IN5VC@?IR*BJ*SGDIR8QYFB4+09:;^9EG>1VD9V-T 
@JC4MB3^#"B=<@%[]R<,-3.T'@W()PCB Q><S]#+GT_T 
@>J5,%=AUQ%OLV'GF*/XN_:Y.#IL_LR$QLIG%W9,T>-  
@\**7V^[N,/B6G8:G9&>266L\C^J2K?I,@"4!.Q#$V@, 
@IB)[@)[4+)#QR4$?^T(5GIVS$;/./MNQM01LF 0CZ_0 
@7<S_#)4,[4=O5_O=$R(ES-8&G/DTW[ZES-6\CZN>K<< 
@><A2^SB'+OF9PF5P[/<F(%W_MA=$)H*7=.RJ7#BWN6L 
@2O SNQH,70THM'FZ#*0IW":'+] 67EH'*K45$R+I<.\ 
@?*B[( X$^^R(_2W7\<[0<Z"HAU-RBH*;R^U8/+!!$^  
@HT9.Y>KV0CQ,(@%U_;(M:&0H&>3B37 .2-$#>QK2:RH 
@Q546[G[D$&^.4P+IJ2:9M\EEZTF[-<&F(CD:8C5ELC( 
@7@U[14$U\9UMU&CELV88D.<X4SFP4TP=GO_DS+Q%<D4 
@+] (I[*BD^]+B'Z:\V0F&&1$*J&(WW;TTS$1N&KIS7< 
@VG7ZB^8#^Z[Q0SO4WO;P&_=,<4CY\T?1"=I2<FY3_<L 
@98*NF_^((I?KQ6I=JRO07OGMDV;-EX898.DEPFQBZ/D 
@3R,]OD.2$_,(U,2H?$V^IRR.5P\VH&&N,<NZR& _$S4 
@%\#AX4QV^>0U2(3V;>Y7A><$"34\>(.]Q@VLZ(>/_1( 
@&X_I#W'K[7RTDM@; -TFNOE6E!9HJ&8*&_24UB!\M'@ 
@3[H?O]O>,R*=JQQR7ER%K[MKV_JYTPJ BN#3D2X$)^< 
@OV+]:&_+<^^.>PVO/$X2P]M"KCQOR>(B1H]N.=_]F\T 
@LMUV\OP;SBSB3H<UR%14+)@B.AU!9(IF?B?(LS38M/  
@,-FNYV\C>$'&6;FU>]YZ'2<M[1\5=SSX=-=U8&K#65X 
@]"< ]MF8(RHD2%XZ/3/E>*,T>'!;4@L _0LV\#1GN<X 
@ZW$@G])DB%JC<_32/2+6W)&N3#')&PX2B6]C2A*O,]P 
@DVI];>NLYF6=1D(5"&8X$K:B7 G:3V1Z*T]\S!PAJJH 
@\0!6-Q?1_C_/I A9\_QZQ<@KF!M[%SXQ"L#2Q]XL'J4 
@(5D!HA3W9I)AU;570+'IW?G[M-/@%$@@O2S6E"ICMF, 
@PA:!V_._?%9N3*Y?-Y^K]]*==XP8531.4-4 D\?C"8, 
@^&EI..=)O' 3\?G=Z2#@1/NJPW-UA34+\6H_=)P8QQ0 
@LBPVI.!_9%CA)0_44, $F)F"_^DI04MUVCGY>]FBY00 
@H^7,_U1\[05_T.(:8[=:+5#EU_<1_&B#NJRP3YAC\OT 
@:5%BB0;*X1R!)R]@;R#Q!HXIVS/LH/[.R%S%<#5G"K\ 
@[^!9Z3@5 *4!H,F:)&:0(A@ 5PK*N]->'^H!U&H@>?X 
@51<LIL^V1EA,O<@6&T$W<$JMPA35R9CH>B$(L#+>XT4 
@QM4#.([/?!*\D4:D:%LFU_UO.6)C!.7U$E*100<YR]4 
@G\OO?"Q(6NG:\;=^$$K$+ Z,=IBUWSXFSXVD:@>3IUP 
@W@Y!=)<L8]L]+"IMKK+"@X3#,W\$/#?JYI"'9T3-5>@ 
@V+:@(@Y2+7>,D?EV0 &0_?%,?9G[2URD>]VB/X7%HB4 
@GN\9:O.:N5HIIVE-*72XJN=)_^_-GK<#*;IT4_4I =( 
@>Q=6_#$J=H;"L^KEP4NFHGEBZ+"QRY=;Z""R7.^$L-0 
@W4S4&V0'1?U)3)H1I$B) ,(LESGL(#1\-MMX 'PWY 8 
@?0/%)H R8EEHOV.M=[U.PY,(J8+ ^M].J%^#RNS*F98 
@&HZ1A/R\Q;::Q=RG\ 0GZ=<-[,5!K7[^J2&Z*:/]+0D 
@O^D>C[,FXM+8?P/=;4$)HKP8&V?]UR0+SE(+"8;S4(4 
@G1(J^7IM"L=)5.8>[L^N)Y'+EK^B)%095L!.\$H:S8( 
@M4[.*^PLFEQ$!HR/N;?[K%&DYS%ED-SW1GHDU<GI^H4 
@>WPRT2JVR0YA5&YJURO.AP'(?MH?*#<1G=C'^5GP7[  
@A[N1!<T1NW#Q2XLRNEF9PRC7_Y/6T"<.9%,3'/ZFZFL 
@(C.^;<D\0?D<@ WW90'[=[)1DTS"=>41%VM+L;!^0H  
@A7?@G^*,*5^S:-NCAUI,[SO=,/0#?9:/L4OX5_.XDOX 
@\N3\[%6=>'Z,=&.<0G6&N(DRQ=I*&"%^U"99,6Y^8-L 
@98__*W3?HENB]]%T=S_$2^UYKLYZY,:/E__#*:VXKVT 
@UB?PQ%P:-N5<+S'PG>691R+9YF*E1L/\5WEU>MC\"PX 
@'#Y<D(&Q9U0L?5@B"3EHZR;<$"M_]<T@5]#Y (F!=>  
@$R8]-0T?++P:0=3X'K1LOZZ,+=#Q2C<!+F'K^=9+1.X 
@$+D'^7423:TV07J\U-9M5[NP%LR#2\0@!-$:\QWIZS\ 
@/;#)@ "G.>(#_B"=AMEM&UYK[8PR4A=&[$-L"&,-3<X 
@(=;:;MS\Z(QPTUKV%&HF+7QTK23XA.;FK4)5BO*4;*T 
@'-QW'MIP!!F!U7#:HB]7\NLV,$!$OP#V658$MZ4K&?D 
@AB_Z$O?$UW9I*4662$KEP]#X]<:_\OG1WC+86>.. 60 
@\6K)_C/P:$YCI,>YX)T)?]U<[$0Y_[(G%PO$KE+/ <T 
@(22VQ23):LYBC7.5$G)+S51G).._P )I\Y8?4%V+TJ, 
@VYRSUAG .&\,.1B'B60<B_IO!&&I[GBA!3Q=L7H:;?T 
@;6=#K."-0ZEYP96'=5/2V*IAHR:RT8:;M"/4("<H7H\ 
@%T)C('#^S#?VZJU0C">/)+/6PZEZ:$.ICXQ18R;PFSH 
@FQ+N&XTR1'^J,V#VT%^OIHDU:[H)LRJ>,(/8+A^;_H0 
@^VOC[SUO:;,*<S X9. V/<$6+F#Z,]'Z&8':IM2CN6X 
@1 ,&&9")IZ4YF)4?K'<[#A0T!:.5&LE@WT.O\3,:;,P 
@#WT:KH$O>'W!K%YOTB3%[%G25A31D_]!1O:Y6%YB?8H 
@AEZNWJRX5+7*LJRAO[YLC'!T@KK,%#@X2$3#9>@- 1< 
@6(KR#/;M)A#88KS&\LZ*71V><]/E,RM:J)S(;:HB7:, 
@WRM,$$7X9['RCBV&/YX.?P [U]WM43+Z;-%R"UKDB*L 
@,3/2+BE2&[EG8XNU92\-A]00,==+$DQ6M.&!OFL&]2T 
@>=T.J<R/"#5< DA.M @Y@S8;.P_^B( H75SHUJ9\53, 
@2^7R<F&+T#G]4\R=I]C6>K(MXRV&CZ0GL3O,[LXMT$P 
@SR8$IR."QFTPOI3)^P#X@T0RYDKDFI+84.MXL@:(I!D 
@L[92JQMO)$V9&XI9K5=VSAT?8FL6!<-;E-EV^2HA+\< 
@2,*G9A))XTPJ&X,$Q9NWPKT4AWJ$WN] I1,!Q_JUS@0 
@)9-?P6#ZTRV1QRAG>G_2S;%SH"9U&/<MTR")#]A#H/( 
@19-[[:P3*N%=RID_9LGLP7IKG1?SIA96YT=F:6T5N*D 
@I7:>%*"@=MH?N-K>E2%.06LCI3GLY'\PH4POITE)_;$ 
@H;I@^JY.YEGNE/R736&.4Q&1W^;$D6\]#J&CL5.)L"( 
@9MCO2>]$OLZVF.2-.3#$,VB /-*A47%Q?(1*DB]XI*( 
@V-G]7(C <^?<P+KI.%O270T^46B5>6<EJ89GE!5[R(@ 
@87P?2L:OXS37#\Q 5D)#M**H/F11M4HX#')UVMO Y7P 
@U(Q:>JOA05OX^"R6(CMGZ=*NQSLD/=B&- >,V+N:R"D 
@Q F_WU[IZ;NUR64*BWD 9=A\X>&-/#)\-+:P6V2%T\$ 
@^Z!!M/XC0^"A;:)YPD?PEC#.W*3ASM3TQOS>W5_H:*( 
@Y]O.\_$G2ATB9;_F=0X62V\%GFAXRHCUK?/J#&3Q9:$ 
@I.'RQ3U6DIO,E2VA>S[Q+.MES9&12!#*BK&S]<K4R[, 
@>&^SBF1L@\5U6"0V-BY:LKI$'@)*-,E6E7S'DRW>C,\ 
@3O'*=*5B5GEKE'[!:++RMQ_I&6_.?\$6O($ R2'=L^X 
@ASJIH,_\:QK\CSC4M5/#( 50(> ]%O;)1ZS2*GU)A(4 
@JVR>'+DAI1Y33,QC$7R2+][V?1GAWC;,V]KLWF/T"3\ 
@/WJG#ZZI<%MH&K:>0]RDS9,;LI7@RNR]N\760NB.VUX 
@?,=+"T3A?MON9=O -C,=G_>96!KUNB1S:*BH?^2SC(H 
@@D6C]FH*F<5AVR7#E8;LIQ7IJ!\#F]*)=1\9;$" U/X 
@[!NTDPK-\ [S7(B@78-9I]&DUN!0U[8$LFKCN>?@[4H 
@'X5#<+LTWNVWFW)?O%RK_&->HN4VL;")^G31$ >#80$ 
@&E$#)*.T#OTJV(QN@GDB,R62[.G4RJ9ND-5^'F:Y*I@ 
@.L1M2%U-'O._F3HNA;BXP\<)_ PP-B/',"'1N?]L,@@ 
@?0+K\HI&CD4/$#*Q;&A<E!H;86DU(4Z'1!J GX3:QMX 
@.S0>'?0BQ40<D9@1V_K\4\=8=*R^VUM85:H>-20!T(0 
@G\M:".("_@7QCH26(]-V[9'"51DBP4X<PL-9DU*[24P 
@T@MFFA8E?"4?^YQ;QV"4;L$DH6<S<7R\A65=\L;_8R0 
@%IJ<*,I]]%/N^Q<B<:J@#TNS#1#U#ULFO5*+7K]6EC\ 
@MIQO-XYK[C=K;>'$'=#*_I&<[L6_=9.A%[-"6/4Q!C< 
@PA204&0ZIAM6TZ<5T%[FA9-)_W_>I"=*G,<>%S$(/I@ 
@.6SH.O 29(O]E%#HM* !IC 57#>-V0<XN,MH-APW6Q4 
@\VPN<U11($(LR5INC\-;4+WG<Y/VT)N1P<:HH<[[=W\ 
@?JF,S6,#L+1:&Z$6"K XG]6;RN'Y8GGG-=%AJ?ZL8YH 
@%#8Y8$^@2 MBM[O(WU&,6R]-EV/%]^86Z2=T!''D8[@ 
@,KIQ5</WH=X2G+KF!',YZU5GWW+^2/#Q?8!J#)OU29< 
@DK:V-+.S6!T0E&L,9C9^\^7JS-T3XW!8[V=:V]EHX@X 
@)^==P!5:4Z4QF)8JO,+0RG8KYE/U*PYWU3II3D#50*, 
@4MZ,W#T/_$H=*6:ET=#GQ?$74&!4(VHK9W,S'%_&*(\ 
@O1%\"?=!N22^82TR-!?$"+ 9<@:5?R)U7K\$B?24258 
@IE>QD!L3H(':K>J?"&F@02A7*507WSY'+\1<)MB64S, 
@E.^=(OWCIN!C1[G+Q?G3,B.F2"]0CA_V/ G'@$-;Y+L 
@'>+#,Z/JC"JQ?V^7RTK0Q$+(3H7C?=UIC,,Y[9$HB+\ 
@<Z!C:S-#,5[J\/RBH6%Y$=N:HD<AXW'*EK*K[3V[[U$ 
@NR/H9!B7!ZFAYZ=2WG/#(IY";Z/ZWAPE4JFF"8H [Q\ 
@]5!UMB;&3NI"4VJPWJ[_$T36JUR<96R'@^BK;#R83%X 
@@?5!# RW5;0\'0# <!'5XB*XI2(S=(?1PIWH-[+\ZY$ 
@1@*N7X60K73<W,$3.O<D0*@IR %1,+E*6!W#IX*1S:X 
@ 75928=;@?=D>Y9D83! S,(6H+WVO=KU4Z6XA)@]HGD 
@=4''Z+>?5O<Q04/7MU"@@R#7Y]E<P\=8]O<QOPHF>!L 
@1AU(Y'I"H.KWRW'<&F,4T<B^I F@V2O6W?V0T-0)!,, 
@XB0W42OS3D9#DT"\Y<PW=VR6&T O?KM#)GLVJK#V5W< 
@ ;$0)>CV,Q0]5G'<6$GI;-=<C%?K4 RRT=K=IA.0!TD 
@,&_%ITX6)D>,MIJ$:NESRH<AK$5$[]/DF[AQ;YBKEC@ 
@RSIIE=("F7Q<QT)#1?9*(8,"&<4FS.-%: _E/&\<TK( 
@S&Y+KYO+#H]$HLOL N0_"<=? D(UET:& 8+I?^G7. ( 
@0]I+5 F9_2VKC7;1YZ3C&OI;[6X<9E:OTQ)YF?6B8XH 
@#(!Q&71Y50Y_+U-3X*;)G^HXAD"2,@'04X7HI\\P[]L 
@;I9^1L&D-VC9ETM=BU^8@"UU'S!'U#!5=N%J6]3J,78 
@,4YZ0AYM-F##+XSV@HIL0QX87SP&G4R.JZWAEJY8 ,X 
@?_ZPI8H/+7VBAXU'&%;V9P+A^FM]3^8!QLF%1FP'@I$ 
@3U /7?J0H3[<Q[H<PYT!87][@<>*0@<8!?9'/= SJ:H 
@QI#.0 .UW]J1<Z3^(H8A:HZDJ50G.JN:N4F;97BU#SX 
@PTC\ J_JEV'R[/,X80$JO2/[5I9("6?94&W<NKO'SW$ 
@0=H(N/@$4J<E85*I:*:O*MIF/;>!QWT7>7GUTAZW0KL 
@U,DC)JIZ>E!5()=Z;#+@*NTXT5#!RE&O.=LA,)I_3E@ 
@VD!(M5F)X*#[6CR(M"VUHOG&%]_4M7]I*'VT9)H"K)8 
@\RM?0XA=5VOKRS<7UK2@?=*L&)X7'L&2N9#X6WC,W*( 
@/&Y[S6& X;Q>NAK;.9Z<8FPC^'NI, RNFO)Y54>Y\R4 
@6$>QT$S-9<F5ZL7"YMCB4L+'$WI4V&A'G*G]I\__'^< 
@=BP)%RW*Q*I,$K,,5^EMDDX:Q.1?%LWQO1H6TJ*!WKT 
@(:0OTR\+Y5L&PHY%:B5I"8*<F <WJF&)^1G;@S1R@5P 
@9":B>A2<9IJ4+K9MTS5=?6C2 ^(5FY2?.-"P[(M*%M4 
@F.[<=;?*1 P\\0]D8YLOZG4"W(-D^0A; $)W[A):3.< 
@D(,$=?!T@QK44R%[E2K:X3B JVBQ$<L4^;=Y9%^KG9D 
@1/Y^4\>_'-MG%[.)708B$C@&#G!%J\J$#;JS&.$HVNL 
@1N.C041GL3/\KJQV?FK=TS,"[_0;%PV$AA.'US==2>  
@222F*Y=L"7]M$"6;VZ,UP.,X18.LD845&X9C3S'G\RX 
@W.%5YW:!*&/<J1D>C0Y7RUY*<B/9%J#\7:5.3]!-E?T 
@N-&2\<!9B@N/+CX9%8IVB3GP,&J+4?B9&G&ZF-#U)4( 
@2N&=D&VDI0A/TG7HR'%$9^)?48.!-<M1>:B;([9[!TD 
@88[P0BA4->TTT)U,H30\=UNPKI'5G)$6Q(B1I&ST_WP 
@+,#Z?DDK)^/B+9_4G'S])[N4Z29<O/A\G( U]@XT"8@ 
@GA&"V&%TF^H+^":/RZ ^08)N^  A4Y"9]8>'!:>GGK, 
@8R'Y8J"8@SS@UN$Y%YYOLU?;N(!*-/X&N39NG'G8;U0 
@8HL#-_!'3/,J*.[0: 3\*!>(#+A!MVZH8<=X!KW\+GD 
@"(HBY9;5:2 60RVH1;PW]W8G& _ &LT"5;E7B(J!WYL 
@=:&Z/%RO/;5O53<-MYAG84-\4R;\Q"%_#_-,WP\3'3$ 
@0E#D[N*;+U2YB_ )J9 ,E<)JRC0I)>5/4A>&D,6D#D, 
@MX<^;I>+89TUM3X#5"4S\@L0>-8,N1DO)\+[KMRZSX\ 
@&V4D8-*Q..87:W5S48!RE;L'D934>Y$E^@2EFMF.(OH 
@\V?HX>R T:LJ.-;+?T7.H+T)R3D.\$M1./DK.'W3LY8 
@T?P<LL\#MH?&#N:84$U;QF8E[_[*M4G_P5?(F$AORQ\ 
@X2$CY\=)#:3RMRU@%\"<AH?;Y!NAE1E_1<KSWTJS\'\ 
@-V&")_#M-7@@<D%*OM1DJE&6#".+M/0V]R(,MRYIB^D 
@R6E*R8 H6#/\_!$T*&%$ZLS'6PXG(2W]KF-;2<W99KL 
@P;G"(3N7U2ZB5JS!M;14L,/DI&ND>:)%E6L C7<L014 
@;)Y5QH;NW,XU:"LX)Y$1O;+'K22RSXGBX,!]G^F+U&< 
@W?(4(1IX:GSZ5>@"OD*!9.\#E"K1"]/6O J;U["?SQ< 
@/-B1U"$E^Y195[[Q1&B8[M=UKB5@N)A2,E.EFT P&;4 
@%*5%*'*K7Q../8+2.>79BQ0K+PW$F.^0,-7_PW<KE=( 
@)3V?=*4 %NW>PN@R1?1AY3*S Z:+)^/G3G,;1JY0C!4 
@+C!$K2:F>59?!R!6]I(0'[JF#DL=6X-Q9!QI4Q3(^8< 
@FX%0C),%M8Z\-*:L_8-9D5^[4$O[R\/TN0M'[U,V#XP 
@!-=JNK /;EC+!FVS'LM&#"A*+E7KTF'L65P#PSH(H/$ 
@6?^VN@IIR60K01M$1R"$? A>)V__B>E:#($[^8[-W4, 
@<5#\W0$C&DB!9M5RU:FH=J0K=4-;0,;]PSDTJTM63.L 
@T1K1T:JF/L+4!/-#Z4?4"XU3"^3WH>+.-2)J-2%@D.@ 
@SI$Y]8U3T?Q,G"!G L#F^QQ^)+=@KKH#+VM+5I#!Q.@ 
@2865O;8"0*)UW'$Y7:-DFY&[^(%1YDO!'@)W[ICA1*P 
@R=QT")A_?M>YH.V\>;ZVJSWXNHG(0C]%BI.)]H&[GA, 
@8<F^)IC=]0Z?A=3$WD0'TC'6<B!\(%;=J3GJ5CP,">@ 
@?DN5>#@LS3_GM+S*XP!W@M;XIE<'6,A9UT#&5VAZ,EL 
@,U)+\OAU2(7A*D[=@9!<F\/B":Q:N_C(U,.A$==7B3T 
@<S*6@,1,-=#6&N)<_1$XIT6IZD=\<-(/ AYN#05;X*T 
@!3=Y5L0C%UI2B0L#1V:L0I/3]T/YH&'8X539-/_K1GL 
@EL P^T^XYGKBI#QL>T1%W%G3?-.Y8FLS%>_WQ)[%?'$ 
@AJGXI&,,*(YG%O>-A5\K-M\H^Q5-=@W^RP]@X7'46P  
@#\)K#U\<;;.97.S72F_PFQ?,6QUTL("VPDL5;@\@;U\ 
@,;.0%ZBIY]\EXDLOQ^#*VZXPB8!356CZA7YT?6EWR#\ 
@@6:G3U#H[$]I\YM=U3 N7?GG=AN0*K36&)YF6OA?KC$ 
@[48ZLKTN>"< )8SI+1W@@GZ97MV3IH$8I,L<*#D;L9$ 
@AR?QN%X@I#%I,5565\N4V6;45^"P/@%X_=(9Y<<0TYX 
@4+C4ZU^*#]*4\9.+]H/+I<0*G,+ED$<]52@8@54=!\X 
@Y7.$,  +B%\0:MZ/5;()EK]35@9E^VD"YL98LNVMAS\ 
@#DQ4,&Y+7+ D  I^@V)R5Z* YC%S%5F,G\C/1L60=:D 
@ 0HG']XO,T+OO?B"P$!W@NE5=QR0%,N7^K@K B]X]+4 
@LA O6>>'9M2O=R400D>T^ #4TICGNL#G:K+'@'(Q-L4 
@;3F\6N%7*,?_LR@Z>H,"FO9QPRIIN@ES?$DB(2L%3*( 
@1;VU:V2,G:D< )1\HDT@65E( @/9R4;T?,*#=^WP>[$ 
@6@2@60EDRWJ-CW6V>.(,H-TJ^D^8\\L7A>Y2#S<A=M, 
@SG";=VDU.&3/8O2L-&R1/B[B6 _#FJ#>47+D#&'-^A8 
@Q3@<<-.P/V/H26CV]W*UI= 4S2,)CVU.9KQ/@O! 3\0 
@7&4;CK"'.W<X<EV*OJP&#B,P<33G[$&.X=?#3CWHE-  
@O#L2(MGHASU^#=:V3E9A^[:>#4=>D5:&9"TO3U=,:"P 
@O:7MPD,"TF*RH:(5VXB1B&O1)+ 6(^[W<A>.TBHB"K@ 
@'HHN$N]'D"#H;UU25[3K5,/?7Y3S!6F#>>M>!R-$8R0 
@>T\$^<$(,\CQO5DC&Z!9^+*N;;%G\]&\_+M@+1,-GK$ 
@&V=H>QFNQK7W WQCJ$4O,5X*=4+N[C;L3-H2M5 T=:< 
@(^GE6763)+M7.1+;_(]^UX0_DCNH'P/Q1;/?B)ZO/WX 
@<#@L^T]-X=^TX*FM2B_51@6SOBRCY/1X>>KS6:=GW6( 
@R I)'9T*))E"2B!B:+&@^0H&[3=,RT0:MO.&3,KY&<\ 
@7FB6 K3@4R.5+Z]BI<W43L9#/A!OU&36<>*KEL@M<)L 
@->V#?S63004#RQLZ!==\UZW1E+S>K9"6!5PP8Z,F#'\ 
@VXM$LZ[3V5?SY=:/2YRBDB[CH&>\1U )_G! RSJ(7"X 
@G8S7UZUHA"F0)QU?S*#2:_^O;[#S<H)X&-6P,HX<KF4 
@7+=K>=/"1C.[ $,E*Y^Z [TA"XF$44X'5$COS"A!Y5, 
@V8R4:X#KL7YHG-E95&7 YE5>,VF%4-/<]+Y 6E?WCB4 
@U'7\_2]1Z#>@\J[8?\4PBT# !?])65FJI ZF$^UP)!T 
@I79=6K_;3K)V$$WJ* KB:#UD6OT+!B!^'2>-2K#A\#( 
@?]EHW7T0CQN(XLP1$AGD/!_S/=6;\Y]658'U<?93&!\ 
@0U<20X$!;;[P@*"$[=.=]B<-,\+R0*8$M2E(GH.)PTP 
@]M/MZ;7_!$(\A[\VPE&JM:)QM3>XX 1+5O=H;WN%N$H 
@UP8_RIXJAM,LS..\W4GUW,!5Z<]X[I0 O*$HWAKEP%8 
@T(.1E/YQ>HX/8V=HC?$%(+PFP[+P9D22%=;H+X$3'YX 
@(V88\60*R.A:GZDJ/0>95!&4/(4%?3SN6#R)O.W!]P@ 
@\JB.&)>5XQ]FSA]WB14UX@I47S8?RJ^2O;JY]0EP_L\ 
@^;8AE_;F8Y%<T#V%X.ORHM-2NB\ 5UT9&:G?;53#$O( 
@;6K'HZS^D04)_]YTZ92LQZW&[9H@BC +&$N3%%=J'.P 
@B-+4/G@4Y/X>2"!3L5"V&?-;>6U8?B, H?7+AKDVX%4 
@ZWM58.4245JJ[$R/[?1LZI[73J<JL63/9!M>(R$\+*\ 
@RLK-9T!;HPEW<CA?7.<^?U5:3YV\5>"3R[RX!2JR+RL 
@\H6G-4(7HU"83;=0=*R4 1\RE_ZK2T3%+H.9Z*].ZTP 
@QM'WS&;"NEPNS:YSL.ZFDDINDUPGN-=2"QS=U)I0VA8 
@8\1[@[T8W\.5.N*G4+2P"N;4AUF>\XA"S48&;:&NG+  
@FT =_&IMJ6K1P-QU-I_1B%J"/R+V#%IQ1L?H(/R^W\X 
@6_$]AG&A-;!#I?MTS+M? )M+:]$-OWE<&6[L=,$1<%( 
@?$Q0JM#59E2U?^(,2%#XGSP9X.@,G6G+;:ONPM<*.9L 
@?=JAH$R( ,S,NFF<&!OJ)5^5(Y\)K2AKCI.+7^17O[X 
@$TS_//$+WM'NS6&'*-7$8,S5;ER%8E62@3&[(;Q(5-$ 
@R^81N7@V4LJ4+XD:1P4/6]"DES%"(A[33YIR[I;<Z$< 
@VAEE0X,J]:'34B) ZIC?3?>?2A(5,YW78O26"$T&*N  
@'436:G[V@A#IM%KZ4L",NGCNI>ZP"N2X9K*#L9VN.2D 
@*6O0MG..B 0S([X#E3C5B.%:0 JUF7K>#48/[YU;,ET 
@R(HN3KT7AG:6^>515D$V+F.U/)*QOT.4X#@;<_D*;Z, 
@D%#RQR4O+</T,-@*5&<Z#@_B5IB)J,NESEC/%*B$$-$ 
@XN@*8L4:K\V6PNV&-%^<[%)FG?P4F9]QT2]"Q\PK#X4 
@WUB$G6--3CKDK(6&7/(B_VXOQ/)Y RC%!MSZ,> %,$8 
@HJWO@:&90BS(XW$[Z-MI^[5EMA<,_-!1 0:'ROS<'J\ 
@GN/*N::E9T G/(B59P8;]P>K)PP2@G1% T@# R:!Q>\ 
@*FM?'2F!OA;/() : >"V85:VI$9_CN#4 -6)^XL X1P 
@^)^ IX53ZZ&<@WPCE]4%:4&,MBLX>%Z-K]()&\,@0P, 
@2R]O:B Q_45U"?1+^?3&UUIPF8;$U8'Z/>8HBNA1:PD 
@ &O?DO7* G"?M"6^4$=NC^D 9;351K2>R-RW.-,39_@ 
@LI.2,J41;6/N/$%GQ%N8TQU$_Q)ISV[E<P7KNQ9J.<  
@O&NMG]]Q:)VS,HA#N#XD@39@)P<]K=KN&B"Q*!Q,RB  
@H8[+J0#+RS)R89JZ)DY3HWU9N02?J1@4$]F&"&4-)-( 
@-2+;<%4C2@&A<X;M0%B*![V@CNB/4H2X+ RT%Q^0544 
@C6"6R6CR#!K98!D%S5](N6J)X^#'%B@0S=.%"DF?3_< 
@$84NF$7MQCKL$7W<G9G)#Z3V[)H'3FTV:K8YHXC%$X4 
@]$0!@M!J*4EP 7%3(5C1NT]KCFC)N0SI+)G6M(;W#.X 
@ '"$];OALG!Q,/[]Q7&?&<-?N_0Y<C4\X27MB7W5!?, 
@)NFX/<_JSNCDQ- [3%!7E5<Y!2ZMH]_G\CH3)A?A45L 
@Z3D>N^[Q+MH +IFD._S+2$ZC2K6$'19'^E]VN04$;J4 
@-<4DPT'*#S$9I&V7DM!$L/((W'1M\/]NU=]]W-9)U+P 
@R8A_!0@JT=3D< HKPJ0%%U?6.,07Y!C;E I5NY<[-UP 
@-?13S5GXJ!R)?&,;=!F:K*11 /:/)REKGAM!SV<-'-4 
@GNU=6?8QMJO>JC4UO!. 15XV-<B=L@P%"5S.4/+RPY< 
@"R# 1&]5Z&GYH,?6*NV:1@(T&&9\",2'/#0UHR!9YJ\ 
@$&(ZDX8+8!-9NQVQ-7>/-557] "S".SW<X#(\6!RDTL 
@=N!XZ#QLT[-!OJ%S5S/[YD?>(^T]8 \YB!V^CX _.5, 
@LY6/)<333_?->$8BJM^=Y_+"-LQ6OX7:34OSWS)IM<$ 
@!]?4'=PIAE&=G,,9&=/3MM'O(F$2\SDU.^T"5H88F5, 
@'OGH%C'+C5(/.J::= /=""#A&IHYZ<?-02WC8^HU5FD 
@_/(=TB3,A-C_>UI8/V8?  -.7<"FVOT&HRNMC+TIYG, 
@,&"CC#A!JA8K;@KA&S<_=&#TXI*$UO N(78Y-9MS=A( 
@ZRI^6*_QL^NM.\\O&1GO-T-TTWMH 1.S8C62^<JQ2'8 
@/YST*;$XVRK8'6-JTL25!?H0=Y=)V$?#S<QG+Z#WD2X 
@@=/?#I*:&TA%3VTR$RKM;)U[79L5"?G N&14<3[SO4\ 
@"I/0= 2D$-FCVN6N-*N575PC_<K![<IJE04ENG_*(Q( 
@MA4'0@&K=(YN;P;V)<X^XZPC7[4D]%U[M O-/1PO R$ 
@OX<FR>%\&IN!IB$GWV(\4(WY.CBA#64X^M#LL6>H^4( 
@V3SA=KQ@=!2GZ11WU8AQT',\)@5(J8>GC69Z7.(^U2  
@F('^PW6Q0V* '9OQ8"JQ*['[C'.=SWG[<O=MOB0:@5, 
@3AO"M_-",R=B/=M5TXRNN[:1[3<'B=A3ZXV+=9V\(-H 
@U^4* <E/]:_X9O(7DDFQT9[O:048<>Z\B#P6]W8M\NL 
@<A0=8'(SQ@#!,)2"?+4/CN_%>EF)C^E=:: C6VB$1/, 
@!^,,^>@-=*BQ8CG-O_<P['[Y/(&Y7^\70MD E0]/\%< 
@W)#C6$(CO<H-]^X)NG=%/3T1ESFD2 _.%6T;W<L-,6< 
@R\HU)T:'HF.&WNE8AY3W>GEOA*001X/*<#^)$"F"=\8 
0F@Z*O(P]. DF1*&Q3Z- D   
0%FDRGUI/P#Y3L1MC)&47B@  
`pragma protect end_protected
