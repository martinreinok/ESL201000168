// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
LPglRu2AqWbfy9rfzeQFj116rXlIDSdDtItQrUCDaNW9eEiC+FKh8NBXnYTtPd67
UCadTxcAvzPS0j1ucYmyjtpVJQXiBY7n/Ojx7iE+hbPJXwGnOOtE0C/GSLNnYS7G
twzKMnecGAbIupnBNCjOr/EXPJozNOT7NnERyyVn2up0q2sV6DugXw==
//pragma protect end_key_block
//pragma protect digest_block
0Bip0+hcz9U4G1GVYUltXpAVPQE=
//pragma protect end_digest_block
//pragma protect data_block
H8XycqbWCk7zOgtea07/qS2y1Y9h8cvTLww6vdEKr/RI3CTuOKSdG0A0eKNay25M
R7SMNCBNFbBWEdG2hgE86+Sso5dW8Xflk8F9NwSsJG0WxPmeqGA4E0OdrHLdhv2h
qitQyeA9IrP2IOQVkmZAuqEFWjraR5H+CljObAQ/fsfX91wUHI9WVLAQ9QwGU1h6
8jYdyu04+2XjaqMyCBUigE9UFJACtJpvitKoYdrO87JTtfZ6CZ9Ass2yyYYxTSIK
xGImrMTo7A6HQ8uL4iRswtOacbFLOvvhdV4gjZn8FNJBwsn0+VEovvRXAQxe3saR
iO5pKzUkh+dWJAFGQ4TQZm+/zogNy5VceX/GdZ5PBBBVOFFoDEUtZ+bLWHMEVph0
LQXrLittfLM3OSX+1SqXKVo3PFoqexBZUaZ9JhscDYstRaw5zH4npkgU5MfEUqn1
7G1gqnjiyzfofEVKqMZ6yRac09Uyv3FIMaCS6tgjkko2uwJu2TkazsBVHNs5FgjF
Xmdb2ZvnpKfwbGYxzeRe2biCNro7mryisp0Tc8AotAFQIMmrMoOPq4nFnqV/ffNp
onEiEyscP5Hq+WwNdLSlaOYfhVlYKPpMkQEGR6lNj4HLOQOABwRrMkYrxmkl3dyE
H6O68dqE8Ni414izdEWF6TFCxNiCCtONy7/UjHbXpCuXQbq5NOM8qWdePKZfJtEQ
tdrz3JNtte3UQ2Jmck2w+NAzodS09o1WKVobyP7UBXQwhcwBRxL+iBaeAY2wHsUw
2AGhLO00mFlJNMk03qJyykRX3I9eOlDAzap9o4fnPbXtPUWjxmMnErM3gfikgSnV
/Lzgi0R/zJU2eV61GrDEzlxXGbgfELzJcLKAWdnjiBpjLubUBpYQQ6oEC8xkk9KN
KOKJfB/Mr0Ei4qATCpuM2XuVP/pFKuqMAaqoVUFVHtCoJYNT+TmD5itcT+Ly6Jd/
J7MgrJBvyP7zcJBVixk+gLXIrGD/GXmtH3KEREyM+LXYZZesyZOD4uqNjxAd/9/i
f/m93dmLhO4yNpXRHCX2ksXtf3fkF26eytSosqerK66JNdY/PzAj5lxK7FGnIMp/
VbavUsg4q+2MbZwV7RyWl99Q6njIPi1DmfEASybe8cGklcnGeNfQZvmZ5oztUHL/
sE22eje39hQBlTsxe1IIvuh0iX1csRLpJ84UYYbOHl/80vfTbMluyvQu722zM2hY
4qMN2cSppXrX2oQ6qfh1gbWDRMvSf2SnURmd5O2ZR5+1E1xspGDkvhZvQz/a75eO
XVm2reqh7xafDvBmPhqOgEOaHrnfc8vjyKZhyOqDp4hGlmtCLw1OaBJ1HJdJdmR2
vhpy3+pfDt0Km7+GeUQudlQRKmplTVGTbd6jhbr57qef/HZ4nNdMRzZzzhNhARhs
oo/mpO3DqcwExF+6dtrsjMURJ9Wum/u7nx3oM9LzfnT+cEWMd8t88VlrkPPNKeXv
62dhDkKMwBbAfAA2QNaLHT7supyW5/Q5D/8rOmz6yBAiqPPP0vLt/3xGqS4gV73l
NIlYCn5VTeSFQzI74IMXWR5R82Hp1J2+10cEO5pNwmNSCKj0QoCvwFMetq5PnAWG
k2Bwz5+M6G9ppY8RkYV0I5IXUQFmFaMrimJhVgeAc7InV7Sf5S93hrkrSqd1V8dD
4JwSjuoDmMSUFsiJtnxv6UiJNy/ltZK8e7iuMSwyNHRtTBEJ5F2awbCTjan71KV7
FJi0uu1NeL6ffx88rGDGvxo6UfjsyQ+4fyJUVtp4jGNOWj02mIHNexc62l+Qwbw3
3shd36FkcSQc5h8AObn51qPT+maoEfqZs+D6ivUMQmL84x7oXOFYdM+tyZG9NOkZ
LaI/GuYMgI/BsF+xgKVHIYidgqE6zxMUDpLyeHwDEJiXsPMMPKnkF0iQh6iFN2K+
yhUnPQGSjQmIw0H1zNx4Bbiez0PDgKzD4E4aMDtiqwDfFV2m8ucERuk+p50p2C5l
JViT8+i8pQienNuHDy3SAnU+bdsCeZzSKF68HMbymslmbm15KeJpJNMQIgA78yry
go8GjTWoOZSyNCmQ4cB6Na3bRQTIzJOfwONJ/L5fFsMEZekhfj1v/r9I0XpH5mgy
1lOW0RIqmdxDkjUbxn/Wc0tagpddo4xUCc7n94RE0MveUvNrPYi1eS94q5tp/1k8
/XDCziE9reZEof0bgGc23pE54Ni9Rut4LgE10Wl0oVtmHezxLuNUwtGK4Ck+jGaT
xLnbkwtq47zhbD7svp9C6Ak/AE6pqZ/QkwZ+IFZSlmQoZHWrdk5hdpeXslMsk5YT
aMpUwvCSjvVi10OrJGBLbk5LFoR2GeEsu0iCKQ4R/EkQxp4jNEJRR6AcRSjoQfUs
HQxq8DsO39aGCgsulfas4+tUzTTtNAwHre+8rWVJk9W5gZblxyZeY9d0z+EvJwIw
pR482lPrnia7gMU7cUU6bx3lAdOT0BXLC5so2uhiumdUSOualM/bW5ytUfLL5grs
aYdLbc0ZY2kUH95HVQ1uNThFLDB/FdrjK4SET3r/K5fInDDVk4P3W+n1BzkYtreM
/w67GoUDe88cxgg6izuQj4ezhHDA16qLK4ftkYflEYSnxq1JtmxqAqV7uZj2sAsD
DABgVmtmNKifsfpWxIREorM0tO06MASS70h+4vDoldtW/pO1tzzVCocVtgl5Nbo6
UPRB8doGX5v5A96Z4E9uv1T5zKQWVNSdPzDp5vzISsj7BU8YvwcvVWZxDYeJwlFz
+hiM7ikihTnkNMHrCj71kFvUWn/ZL0J1Z12FjNEDolQe1CWaqEGCZE7CZA8lhEOM
su5WusOoifLTNqKGvcyoh+hS+rs0x+OlhjsxfYfJcJXGCQz7VOEk1KXoL7Ysk79z
sUfsS9jgclK8tuPmLOEi7fl9bjHWE9Q3cwxCdYHGC42ud5NbdY3hKxzKpHk5YuHG
ujPQ3owKwT504QWfaVQsj1h6U6rIByJ15FvdEctEIEXP7jvPn+PclbD5qXY/PFjc
2Pns0Puw0zbM1CEXjo6SRSVJpRkekaSRhL1nU/+qzAgSHiMuDpNVuCIt2lIlwjqn
kWsVYMfCAH8EiBkHnPKgDG7UuLR7yoHXeZVy0FQFkVKlgMKTzZ8Qe1SHqcfgNkiM
ek5RAz9OkPfFk8Z+5K2pb9/QENyUFF3TLGdNXEP6X5bO7vI/BmT85i2uc67pYeej
V1bpR1+fWnDtOmrvZkzXDvk6zoVsMY821SF/GvRZt2M+8LXpg0ZxV7D7soQnC9pC
zkA28XiIURvxDd3VdU8a95XDwiukYi9Ev1T8wX5ZhxrQXHMCRGjoFi0M2hRaFbcj
RDF5EmWk53TH5ngYLQ+w7kx1Z029jaToGR1hZmMfgn/Humz7S8tSDB8yI/qwj7c7
y/FrsZhz+LJ7omIbiC3qOag8QQB50fyscFNlVt+9oBI2Z6I7NFQ+sGLHuV/k+igV
ZxkdRawJNQrXPyymEIfKbHG2qRHWhBuyCeOocvtiEknq5EOZZR+6+GuyIKaLNl85
aHew6sB+HRBPD9+t2MZpxrChT+B54LnmN4cJ2qvf7qY+c1+1glKrZvMzEsig6g4q
W+mcNwj8XPFloDE2cXgdc3m4Y1ZSCDq01QHLXuBctDbCy6iNyxcsHWVju88GNstb
BHKfr4Km/RNGlskZdBo3UPZ9ZvZH1eLnrvkVoCOUFv7UXnIV80bcYw2Ucpi3lht7
hbXzK+Et1tm2enJcNYAwSwKHLFjkoEFBRPc1rVX+aGPQpSCggO0uwvfgoX/RX00V
yXC0pE9nbwBnbd8KMoONU4tGOeb3ooorsfElfCLpRj8niXwXOr+nTXPKeyUDqnf3
F4rz2wNi/MfSu3MF0MKg6rG8cDrz9faf0k58a3rDWbPumQOK/k1GX/GQQEwtlTCa
s75Gu7EBtRK4IzHzZc1Gv1sOtFtEu2fLSjHh3fNmOGueoCutOBbzF5VTvQjrE1Mw
CLlnoB4dkRKknYQDOota1qNnHFeKR+KnzwpD+PiHF/GiVMxnsmBYBjEngquslMHP
BlpQRxyjeC3eFyXOP15S8tiaDVZk9NfzbPTvGRF76RiUWa1lWtNghu5WIAc/ifEa
nwz7jlOIPZaCaTJKj8O13Wsjl0ri592gSK1okoIXHQ54jWSYFevwj1d/S6+mlNkC
PPsfQYbbd81kYKATY8OMMtSGqxoSmMdabvgA2da0c8OIO1c50pRncRlUOwvEMK0V
QpnIBtZWfn2rWIhSp+d1aaPg9v1NWMDeYCmpcN4eIgQahkIhs6oCM+L+V704fzrX
YPMuOfLSsH8rZeQwL+MXLDRKaSi+aqxWVWgbAVwrvzkLkRgI6WH7BhdYoVSzSZR8
0EvOozHs43pC5pbt/Yvem6KzscK40dLRIwpp6ru5L2lfpQ8xpDQPrIOIZLzi/mhn
ucx4UjuQiknzNVQtkZgjiVaCfNoig2iQnFBauvodY+Ds3xq1GHEMSkNrS4u1N3Kj
zeZ9lpXGvIXH6GcdIXMMJbAiYFbR/0TXEQ6m9t8rllYsa8U7o3M34yFc4k6NFBCT
mLIniC0eq2HBMAQ0B4Au6Uxem86WWZhpEotPunlfpZAIXuh1VNeb44KI4HYBnlBO
nQQca8qOljyhkRbcoMjWpiOdYZzm8rtaUsRKCSQKlOQDaDNaBpvejRJudDrIfHkj
hxXZHFcRxy6HQDlgS1BOCb51wXWYIqQGdkvp5Jd60o4StKN8Qe/1glzC4tEzHEJK
SBj5IHRrAdELiNKJrg7plfSCjaeHH6wijG3XDPHTv+YiV12bcMRG4yK6VkQ/oDt6
CblBZpC0MC79gYiNVJuamlAZOzucpkX7VKg+FaDSGWYibFHAgwRpfNd1TyywuBOH
2IFyYf9YzKTNUYZBxOMD2A4sonFEFp9j07BMpHu/Pt1v6UTIwZFvDHhcRHp5778v
X5/Zn5x78AUaoq9+u1L4wLmiXnTgHkf4KsNcyOOH86M1EbamOKEOgrlEGygGEBfb
l/TNhxsibAeim0DVasFMFjiDPeSEyCGfMV2yBURvcguLZLZXXeVO2oQ04S9yyOM2
ygbIXvPP/90y3FLzwwUVYtlx06uMJ69Xe9YRaQBCmtDYVMVlqngZcrqZoxOc2ebK
c/J8GF4x73hVHbb3/+DLk6AI+ufLeDrDSerE5R0XqEpk0/5SIqUgMaHECRNO1MQF
207+VR1pfwCOBZuPT8oVoZ8g+c1V1l7wF95lKjDr0kAnO6hdhLZxaS92TkscyH0j
dMuFHKj3D4YiIRuyEFNfzXZ0aN72RFbTFd7xZZLoIMsooLYJUlbjKbBZIRAcdjvX
k6hQjykIYTavnL+VHACjZ4GLmnSRUrisnY7b6Eqcips4Q8nqEHtbugicTrsKrGRJ
6zKcAdwUxTzX0Mrxkf6HUDsF3fwBi7qS81m9y8xt0k4iHF3aplaeeSS0n125JMX1
Mad5UD09LWRYO7YtTXkBm01Y1KXCjkKcVFOZpXLRHt0TPuddMkggOqbUKay4SLWr
2na5BByK1JGgUZIh/P2NobtIQurcRgg+hvsrjKzuLBPk6foU3j5k+eGRJVIeBk3i
yYYSkqTA7hyhPBvZLmITT9kzVh6FZwEMTGPY/jwJqZhihHSgZcqF5nV3iZtobIw5
Cs7FiCAh2u+lTBcqwGD+mrUa4jakCvb2vG8UfMJshehb5bq6PHhQ27lkGu8/Y4RY
rh0gcHToBpfNKXYhiV8qiJVEUQYWTlexXW+/nDlMhdEbWRH6PO3B9UBlReJHcNg8
xE/eAizxgYIgHIBBG4HAEqMOt/usrsj6NXCiQ2j8pF6VysI//faulINSRYp7yt4u
Q3/QA9b0xtYkCE8wWnNKUM5tO4XQ1T7StOtLx8SzeMASSZf4veQoO7iX2NRk87H6
wLWOIDvjNE7TqPt6KGx+KD+kT2t98zwIp5hyybA3fQ1+x1Vr10poeI3SYoABbUyq
GRNNExM5h0HUYad+/cAIRWvXZswoM7GnMBHu1vdz6hnbWWYcf0Xsp47VFlyXRf+U
6MKv9T84VShX9lgmpIQOOLQH9IFXdWnWUKSMnWkGS9Ki6gCNW334a9vpq8wCLVnf
BHV73PSLFPBiOTWr1jv19gZsruuJ6U5wBmEKqhrtZf7FOz63e4MsbD931xqpBtiU
C/VYVtMYh1d8R4lT5p0bjoKuKqqjU5SYzNqbQ6Pf1hZK/DY95QQa4kuPSZa6++0X
eZQsI9IE6oYtknOWVWg302+K0nFXLKEfqaoRTJrncq+lZrfZPFvhOPdViVz1bu65
PHKJLXCgra9YlVeDbbkBJkSsWdIdK3QvDMN/YwWWWCM0upyNoju0XBt8PFkUgVuj
OU0vVF9HvsIY8FgkFJdwbrCPRIHs0/xTi4OLIDhYSXTnLYIADsffn1sGmostoIRC
cIZkk+Go5VplL86lFv5ZV50FWBLdWnO2tIvukj3ZFkm/YHFN54ulaa5JpQRwxBJ7
4FipiYDCpTOU6tbBq7iYOh+xYbb6l0MQRyFUrEEAvM+I9QJasCnM+aOz799+M7SA
8bykVQXAUXe5W9b7tvaFGQzAFI/gjbNwCxk/8KQaFI5LaLwwVMISU7aYMcJLsgrA
F5HNShJd+zwD4R7qO89AAnt9SnOJCX54B3i9pJZbVCkDCHQ8zaE9GGvvBeVkBL8M
cHMutKA5Y1hobuF0cuagfbf6xXO2+xbJTFgS9TRmhBtY97O5gSVjIGYJwk5Jg1wG
pxdIiQH9emQUQ/HNTnJ22/3i/vJJm1x4GeSj/ymOD8PVWGimUFCD4tRW0YWSeX8o
EMeDkswKd7l+Zdlk4B8ZGRYmFo2uSqA1JNLL8dinfXe6r85rlmAsQxhaP5vyHEKP
TxDlFJZkJd9k1Dm7m0/qx0mdg+GQ+GPS96aAf95EUitO6VXbMRBa4BQKw060D2nY
bUg5QzI7o2U8FzHafa4MpcGDuEoOH9BeN9+la8dc9Ps5jS3mxTfjXm2TBdxUmsR/
puNv/RyhVOj6alPtk1h3YSXH+2o4IAjtmz6Ozt/75RngMZ7JfFeghzzL42bVT16Q
DdvqeJu4Kkn1rbkO5qu3M8DmprSR0VadvZCzSD46PLZep12yc4p5GMU/al4X33Ix
X3e9nU8DmnmMswQdL2Loij+pWpRPtXJb6yZ59cfqgKndTjrAaRwlihdI8A10WpSK
ZNAyRfkjAgCb9cImyMtLPeEWtxnomag3oBdAjCeIiiFs52LMWdjk2X+BTrfsDqxb
kKcWWdznUTj2kcdsy89makzQZxNnlXCeHEoLki//GRagzy3mnP3MInoacxbN7k5G
Q2IV60DCqjEZ8D71A2ZTsvHIn+3HsM1qQldAOGsleFj9exhfp94ZThSWXnxQfLvA
/E4FZ+ImGoeka0I59aCU1f4G7RV6ejCIaxvtlMoWOto3VXP6j4evkbhqX4px6cpA
QsnXkFnJaCoVmBG2TWDn41BsStre0/mOphIRzraAT26qkwVIfTzYU5TOrwTlZr24
chTNPLJcG96PUENU/h1k3wGW9EL3J1rXLKS0gsomwF3WG0P7Ybw5Mci7x1MT4LB7
emqqxO4Inp7OGreKgRmm118TBZiV3S00jlss7/nDwLPvFJxjUKK8GAX3/GbQNmeQ
Hcbjwj+Q2vTfBXFK0Hy5ETLaAKtuOAv5f9vyo4Qb1I2gbNs4ssgOxNlr0PQwjxeZ
EvgMNx4EWiVXHngN1Pa7qt96auy6k8piFXva2dzpBBio9AiH3zwiNePnmGpi/pDa
qTVuuz2r/DjCHJob+SrY2bzUK8c0VFJZ/FQbgOnMvem2sVow7Sebm0EyGOXX9J9C
393j2Ba8m5WfzndgroVKss7CP+G04Fh/DTjCIME4I00FOU5T/xgmJXPjJw6HdyDN
k3bTyfwro6ETI0RKPz7NmsJthnSWq3HnQx9x3dKYHi/PjfbkNZpwSN8uvJOT0yQc
Q2Jhrg0aSVhbpGHPrDv0gX/8rq53EtCHuUSgMPOO05NnNIU5rZXlSXgZbPYloY8v
imixAW85O/Tm/+HYwcJ74JZxZGVVsa9Tu0XpECwVezo54eWfyT+YIcmWQze3pnDr
+00455i050KTe8Tv4d4uG+CgF1JkKRo7I4KGGLBup6U+4KMU1zliseavdXEN8ZAc
lojuCxiC/rlztJp7rUBWZrV2UNWoV4CT+Slv/7xRPwZvFdd02sdGEclqVV3/Aq0a
iVctDuT5tWu3A0zpRrqC7RESK3LlJoN90y1VjIa4dcjKb/Od06Oo9V9fXZa2LciH
Xx8eL4mZ6PkqGC7+nJCjQYdJJ1CYc7tDzTK/GdeegIE2otbIIM2tUjFwdh+Q120k
Zipn2GBdYIy9i/cCCOT7v4+Kj4RQi0ghzcohwiSlv2ZkZw0Gepp3u3gVZti9tIza
uwaarQf3Qz1A33XFcLvWtVJBLIN4QPzkKmBfIbed1Yt9vn8sAQciki4H0MXMhdsy
uEtyEZH0qyM/iolDSLxQ2w8nmO10u8yfNvvA+rsSIDC+DBIaeba/Fvk41gbVD7Jo
XoYcMTpPdoBdHZhbnaUYOe4e4USZ69YVTlFx1e1z+8zlApCMJsTV+DtKcWwmHUdd
XZG+GdvK0is5fStb7HOGjCs2BVUjaAfKiKTc3n66qtyK0mTOMRRUeq92CN4Tpd8n
wwvCeXaD6zJvPASJfX50ubyoeT+bvletRvDVlTwfxF3L/N0KMR8U7XYWtX0YR3x+
FT+/iE8kEiL+ZjsCqFr0QWd5pyS8A01F/bY4KJsYm2UCggmRBtGfVNpsqR1+2S53
QNMpnNkVOi3wWujeWxmQ8gWJXhfWhAOArtGH7Igs5YkNXZ3VOaYWaIxCWLAeMhy5
M1Gx6LGIF6LYy+IXN03QTGd9KqFGL+65JNwWBXyCXMQ2L5dpzM4O4svhEbiuEhaa
oRWNaxq8sZJInoIuYmU2GXAJXRL4G5KXstpti+jI6rXcViJv3ryDdUtXwa5AimwA
w1n0Js3iEwIp8es9+/Y+4lMwGwdYsWqa3GfgY6zOyRwuA739XSaAIb+j2h3/vSmK
fFQNGRIo1VaXslZ9uonNJXIgFYqHZgA3QhTYiM3s/ITVnb2WXBlIoCecmjl7mGGk
Lv1IJ/r6vrCnC+QElqz6wPU+y+Ru8wPeqhVJtm5xLmu6M338NSgFklRVvkxZOKmF
iWl2Cmlwu9cDoOS6bhdwUTQGM/SKsSuGViPjylrLCDOYIZbCYvr/OWQyZdrmka8H
ji4c4pLQNRCVRHLi/VLsZlkiZgPk/klDgou2JfWTU5N+AyyKuqctgP8mPUm7Ujss
i5LYxa7nLcox8p6p46oqv/LrWwkaS+TSN2t2Vo5GsRUyuU+6fbRDJfxQiRmQUJj/
K1Goldi5gx+yHg9gVMnTauVuQ0y04ZfNKBw0aR5KwiBWbRe2lpjRQWA2vt5WnC8+
qbUKZNUMcfepuO9BlYC4WgAnNyP0n9t1mOCvXYu+HYvo++ZepdzPyZeEFafOrl9Z
DDUv9le8SSwJJFNEY9c5K2Z20wP9qNCVuwJYbeL5YLe9tRStkGfl4mMmvu6dM8cV
uve6I2Kpq3vyVeq2xiuYUvfR2gyb9WOZo7QtL6XddOdn4kY9LLyZAsWCQWCut9bP
cPFEE/WteXtjEzeCiPtWfMtvsGhjR43ePejgTAzAHTqxj0lYnqSW7hHD1mG8mFXp
tOq99T12FMxismo+T8S12ukJ5NPF3P9uCT01vEtF0g9yjPpH4EPsc0ujfmgUW2f8
foA75foIJhdTisuio0yWbK6wRCoaHJ3f/DjM85H/BOla5qq0jpjnAa8xDTvuoOn1
2Igv/J712SNtav3Q33Y54rEqiyPnUg4ibF8WM1vVoDzFOvMvW9+LohGxcaExKydp
l94LDYYvl+xQLK083mDIfNAq9n/WnvVQzky10wgOJwj1vgQ1Zwupgf1mAOB/0uAv
WJdY9IbMNBk1c/mYZgVn3533us9UtJabyfdHHOdLHL4UeOt4gxbif1zX8gCyXjCR
24OFDDIUWA4ESTG/3T/LDP77paWQr4VqeS0QoN8slh6IDJjAEiZHeCuIKacaFm3c
hCixwb6cO2qwqn4HUhbE3FVKkij90Qnul7h4rS9+1Harfl7DrtdgR/o5XqvTrNTj
MBCKIAPTwlql5Dimg4WExpbRA4+ecRXv2XecrsPxM69WjcJmNKGiEas6Ogfw+xHa
BrNU2jVYW+Qz2NWcWRSZg2fXoZDuN84qxWHf9IO1kT78ajUBtKsb6CCmDdxMDlVr
orLst3+M6zWfITGpnIM6+q92hP8/AOiJSQcA9jHmeYVuub471XZJVHqzxVfYxtHc
hhW5elUrAaZLw9omEEaGcNWgBRqOSo8Ki+S250IzB3wu0HwcnUxlcvBwO3D82AyX
xIQP9+9aBzxLvlMEHBRA7nu1P9yXaEO3L1DqbN/6TASsqkh3s+e9GUEnVgM8WcYI
ZNfRVH84nwHf9BZsMVtJdJXGpvpDnGzF3yipBNd0hpXnBtB13iobfevL9tJBPIO2
L61qjbBSFa7G10/4UBMeiy+Wc4ESHUOV8u2OHFxN6WOlBzIrvgN89kau/yB/6Gkb
XGUzsueh6H58oNyYndT+xHSAnLkiWaetCWU/1ErhPXPp1aYxhAc8MLQ69tk5qBhY
WF2cHG0h+w64o4eLYyD8h9c7d/+twUPRlFDozbfU8TJq1mN/ecxET6zKD8y78ZvT
cXOZQ+2abdseO6QQ2A8NCpbW8vZp0pROPi3GxxbxotxknqBApE4JHeQkCvksdTlP
jGUTnhLrMJo/yOXewJm1UK6VaafKQ1GsfdDaoGUnzvToFKEtf7M0R9+rDHjb5mXi
WP41kzRgNaa7MVbaiRGOP0mqxGuBdZc2nB/h8ngoBfZJmIzJOl/k7RUp3vOSAfUJ
HXanaqeF3Xnmn+0sder8NOYgTSY10niDGiLplN5YkIUbt+pVxeovoE+t+HupV6y+
MQQe3ergMwY92itftMx720QTcfTOl5pFmQFHeGk4Jm0NME9ooNX3Es/RhobG3jEQ
NcIOK/uG0NUEfL7gvSCr1S7pjuRUvQ5gNRljxv1wrQpwzt3zH4fGrK4shYgy7S3p
1Ee2wdOKZnjrKMWfpdGMqPPRfMBO5AkqpUwr24ar+JFdZZwtEeNUBAuGGzTW9DQC
Z7ZN2fymg3nJlkvOfOM6BG8bcTJfiqRioQoVjU5oy0uvf6Ux7RTgvY+d7tQHNk0x
AGhiqvf1OsV1MC3EswQa1gjaxnbDRlzZfUIB9WsMi7Q7MNEH0ejPlR990WvuN7AS
xczQOkhfIuWjNQLy0yGZMHONBG3xcyvxPxlNjjUDcUZU97/0WJRY2uSX83CyznXY
bzqc7sFcVmk8BkYdd5qolYYXZE1WLHMXiLbu3iCB7mERZTT68NWPB80PJjvYE+Vk
wwrdtFcigCczz9Z1K9a0y/LkRjD09CP10B3+GNjy8KZuaZni5QcxsfYGIehbha1d
FRnGmcT0FpdjVufAXqAP8gbnsAvlA8ssjXG857hxXCQlcAkHnuuxk+uaPG0bZrQh
BPDqdLn4d4uHAC1VkNpuLwo2eafiTRtI/Iufjl7iI8gJJACu8c/l9PzCPUNY24rN
1Z0dvRgf2UGku4s6vZ0xNliFE86qck6owL9Qj5uoI4zLvwO3bV/Daot66HZo5l8k
hmFwFIkyPL5N5jCZQJefK2XJI0SzuWC3XAjGdfEoZKHHomGlCxj1Vfx5hZakyZKP
/JVwSGWF6foYpnsFjAr/1Txo1NvXhq2dz6CtxOlXRpE8iMOTBb8PAVeni1tV2cAy
byybfMa39CHWlGYVn8CxAqCUMlhYI5hZIahTS+ji/MP6BORNsMDqFxGaPpnuk83k
bk8Y28Mfd5Lc7CXc9NeRdPkBpqsxT7uFKTa8cmfBLaGcIeSLonWWlXFgmVE1X0o0
aaGGVQmZ4+Lz+ccG+o4wn+RJMwWuRuFZFgpQ7BFx3SvPp0jXjDfPqBzlsTiAXOtw
vsvbjyLHZ/U2F71op5Wwj7TUWvWeXJMV4IkXpgV48ZN+4aCNY0A2n/8bj1l75kjo
HZvsCAs2VE6aUdH4YgC0eO96fPPfvNvSPUJAnFNL4iT9twa/RK8ZQ1s1jB9sZoLy
6YBpytMNGF/o/AJvpJFB+AR6V4fFCRKAwSrK8tNUfJKUrirwdUGw2SGd5WjqZM7D
O/JA3pjSmOmqHRprnpcYhcUgAwNdZKSlnanTcZHfSOXf5ulp0KjH09MB7Uq1XL45
LFZJZxeURcFoT1lFFzsTAy+KDSNfU67vcRpBQf1HoQm3JSseQSf71E/p9pXpRXEd
rj/avBIt8W5MDNJHUFicU9JlkTp8eVu7pwEtjweme++NeNEKWvvfRPWIJhMxh6Yk
qvnqF8coA80uYQ+F5lkPxba9/t328F1DaB0y6IyGcnSc4BgI0IQf1keEDG/7wUb9
1ndSCO0ebQY1NRl/yE0Vifd5v5sreQ8e9fk6bFOdHt0XrHfm7FBlaxFTzm9cIJXW
b6XwdjYX4fdF6hrExYfvZkCC8IUsl/wGmbdbUVfUeZVldytSDodXdpIyA8y2Cmq9
ZwBnkgXUJFyXpg4y3jFBWz+AuFLX6B8U4FMN9/lL0PTtlfVp/GHI3oYGSWCMYhUk
IsqUWbovDbLgbbKdxNj3Su7/xxRLIa68fdpOcoj/Hv3cyL0K1UQUJHEKSWfkCLeo
cRJQTk2AQejGMV2rH8MRmxlSHiYV2qkQYtpo7AI8nCchUxSzyc5lKNOF2l4jEfr1
Hz9UTjTG+gWeE+tdYS5Ma/Vdqd+aM5rnkVSJIszqFrDMLtpg+4deb/PSBYy2RrbT
AwUsr7fcuugGtkz9nmM2r/Rc7kNSGAe1/TiRebe4DyxhcAFHZ7Ax+QzOy56vCRiv
oawe+pdRAYTwvdk2Ktt+bhvMko3PCZBj7JkKlovlF2utnPNN/sslGT6qxCmQ5MzH
FGZoAdjQu1bqrLAruz+9cP/bhmjDByQp3XRmtuErrrn4xrD0C+XUskUzrt99aJgu
N9Uu+7jg3Iw5hMF6i5JP5ReURhHb2NOGJ3CcnMZHiZwnGZPBmuT5Q+5m+4TauQLc
l9jRim1ugoQ2imn483FTHrnG0ep0xtOtqCwThUdPTRATFFEsfCNLa+hhrTlOX09e
Pdoh+3Ca/cUSoOkVW3dIwS7GEMu3LhdQX6Ps8YAx5arSWu7FfsT0JX559kQvQwF0
SU8qHUqIGWOhXOeueqY1+eatT4Sq0TvticIcqP9YZVgGq4XUnBOTsBwkuJXFwjaP
Sd2M5GTtHBrLjsUe5LQiFntmcNM28biELafiXL77sJvFWq88WWKgBupMZWdlXP2f
zUz2Cb+xhCmlTmLpNRas4IinRq4H+1whyHXI5BL3CA2V4DWMT2SrXtTcy6/QmCo0
IRp88ZGwB1a0Dc1xcVL99SKYOogEDRST24PLj25MUuZ1SS8dZwpBtMebS6bKY5eY
Ri7kQlUfn/U1GQz4KhRZ3DFbE0aKi6ACxSOLv8+Yi2V8nK72//Nci7JUMGTFE6CA
CiUnWHRMJUgYT4XPR4LA5NL6uEry4K/+UtX0WxrodQmSijfQRQvcMe05264+tpm2
vDiYUC1ootX9gc3HD7UEX2l1usV2Y+EYymO2icvM5+ZqBaY3Dx1/aq/8ZpFr3SA9
EIZCkj1FcMtBb7lMjjFf8KooezOq1kc2KBVg8lDq0P5I6zDfUqNHloeU0yLs2eAr
jKZTtJ0UNwYTyKut6Mqyaycr9Y4j8XcnMbHHV7GTPOcPtkIiDHXNQ4OBuqcQJlHc
fBXEYGMfhoo4oRLzNFGnAXISjrF7XRV+XrepopAivMoAlFfm+2AgH2QvQSd95RFp
BCNR21xNWa+F7+sGK84F36n+d9yTwDzsUlT7m8JF9kpvN9F1L1+3r8dSNXehs6Pv
xEirLPBzUdw2c8xTf6H5tbvTktNMH7KgYoBeFA8dyhX3CeTmPwowXwcDRrRiDBpw
Whp2q5WYF8ECTEqkB2IRN3iyGcJh2SbdX3RnjKeaBRaGOpRiBaS1RUNfLruUy7JU
Zvu2elLwEMq4fE0sgjSivXgXgkw9wz/iRl32QAIaFZ20Wkp21qIaklhlktKF19RG
4gOY0dlm7Ot3/4PCOJNGeufIe4ZtiVDQtAjeiAqDI+160b4GqfOlajtUhMuZ1Sfa
Q3/rTlEQfWAzZ5svGN/yE2WhV4pzF1uo/0hcaAzVaMsyKMnG366x4n28A3YhK345
Kify+/VtcTP+uCKU2LudY86nwsQuTSQuPo1OaZlT3LRoqCJRfJPYVFezKGBNdirc
aIZyvtnix4X5q4BRqRH2BjUU+A/V1yf9BkbwnkETM8V+dZantu6sqZUMRMwn3liw
ENMCa+W5XI2WKrYdm4B0TmWRTb6waRX0z+EKK7SbIPv1C8rn++dw8uKpQE1PQSrV
pQa8sd5ZAd/IjsNNK7jGL1COt9sG4U7465zCIRY7ie3Qc9E10DjA7RuE88yoQ0La
uY/GiPG/aqaK8Ia+v6qxnRg1jvjhwR2QcRzRlsLF2tC9yZ5tR+VVcZD/KevzKjzR
kBNHWRkKMQSGyRO7QlV50x7TPy0LLqTqbiVxohgB5z3QKKNwbqFOJ77vZrGboLjQ
brRzpLWPAL/UbgeptNpQwp/WKVZ6VIxo7FrBYqIQeJ/Pu+j2ZCRG6h8Ox/YIKUeU
312iUDwTtbNK1ed2kwtB070uN17ygXwgEB0ALwVPiGqOFXrF+WSZacc05i7g337h
5N/It9wzfSy8VBO6ll7rK2hpYcnVZQKbXwBaFiXGm7j+x2i4g0jkLAVu3RzC+3oi
FZFYIr7lth++4nOTQYCGShD4wwfOG+bITSjL2hE3UM0rCcuk3eHn8iV+HU+NYFKx
xmTZQD73Mrbv0LG1c5jE1omi1iZprIneL9FW03Ib3TYCiXY9dggTiDC66BuBC7aS
oDeOIlGtHlY4MekHDB/cFI5igLTG/tiyYgtmSz+mtgnHVZ1ZlmmhlDYRXNSJTGI0
j9O8WtGwTkq6Zshr9ugOvVZ6/yhJSZSPRVYWZD/WPBvnnyAPAyuRCOjx3uwlaxQk
zTQRDZmgefFVUFfJ7LlyIWZAJ/yotw1/K0gvDSmBeBf0pHtwQhvpj+MkgAft3xqb
faPygmOb6w48NiVTz/il3B5D9ZlaCb5K2xH2z51cdQhMf5f4/1sZZxV0Lu41vYps
S6v2kca6JXr1V1D6ZHPuoWkAdN5n5eYHiw2lm3NdMBljDn+cnmIxwda8komfXq+R
mdaOcnr+pZtRbrRiBMKWcBsZq70mWTZ72df7jOzzoBqAdJ6acr7WO614pyZ7QnBd
kP3asOQ2D2KL1Uk0P5TcR4IQpsAkBBFj0YZfRaCGcDT/o0PJZCDg/kR8iH40uoUe
C5SnAIPiMzfgsQnNnhuEegBM85jDwaGIaiO1e78nr71yoYMsiwjtzZTwu7s/r2nP
LHj+hpEvBO7/XaFnWGei7tKB2ovg8hbOpwp0EitFrEpU2Qbh712plpasfvq/3uB5
kjYXA/II3sV6wZBASi/FUCSSIh12IddLQTYTfzCp7ASKWvXloP2yh0Ijdxj874rH
Ni1symL6UaZLrpR34+WLTiK7bGXRCJ4PoKiSFb+BBEHsBBTPMz2b3Zm73Mdr8PwY
BdYppW9dOwlqDz1lnoI1m0jrt/BxB01RZ6u0AFXberytZa+ALk4bLh3nTaVbLRtf
Cs6dP8WhmCP/dGdyPLamYG/Xbclpmv8/4acaiKgGdF8TbIsrIQD4BJ0I0oG2baRI
zYH/8LG8TYJ/TzBpXTTzyxh2BgvwMa93zJEFcpUjkdYd0Asny7fUH8aeDc8QYkpY
U4sYTMfouDzNyonyb+cXvGby5ErlJ9j4HdYTgB043Hl/3ALGMnvoSyMPFq3jCkdc
Hb/CITojbXwZBGu1nG07xQaRicABQpk0ufCDQtYyWfc/KJ7rTJ+zE1DQ2s72TWun
uo6frle9MNIVH2Yp8QwtiY5n94hGTWEDNRBLta3NErqdiYJXbd353/ujenxw+ifE
rJyVQr23i8PmMqO0+BCdFMxIVRdw+W+ePOyx4oxuR3LwADm2cRPseSepUSVEIu56
4YE7FczW0inXbS430znvDoaC+5thCXzPqxAM8EIQ52sLKooiAYmlgl9SMKUVlf4W
Y70yvTVgaSF7smc7lYatwFJ8YV1Znh2Bx4/3aCvF/ON3dw1beKgGaKjVO0Y44aXm
DpUKTSyCvmE9o076xn7DMjiYXFQ+AbilxRSibXqrzGIjr5jGNf4Qw2BuDsYQzRyi
eGH60ODCy7aZRatmUwrGJzaPBU4gKBnOkbvTGEoPFliluEsWHE/Ry3hEbqaSGjU+
oX9zPezLd5kFLA2hlykm2PfwOo2UBk9H3zDEAuLBefgEmk2dHmhZ/WKm06DIRK0c
5QAhf/HODv/1H8Kzkp3Z+81K5S6Wkg/0cjY88YAWiPelTowUL9rXQD9j0cjismeN
m3uszjr0Bd+ohnsmkB+FrcqqaSngPaRBP78ujCK5gR3jwFqeDaj0RqjSfQq0LtMT
ptI2ALIX+tOIffj5okugrCATC5NeX325PbpgcB2x2q++UHe5+01My2USci2ZyGMB
FIgMoMVL98PqB1ODyDdRux8StaxDpGZWg4bXYYHGDAZ6AxvB6an6HaBgfK3CxQBG
S+c4JDPyJZuogsWLjy+is12kK9n5BxD/ZZuIwFGuN9F9wB/SEhXyjBcq9crnvrts
1W855vaod7hnoORIFR2l0FHyHtsjsgtwd/LRMOQB1u1y+sTH2qJ4WqSVybzLH40j
JqwQzuWYB7kl0Ig0elhyvE0yIl0d5tWyUnECVQ+uotndDoTY/Tgz4t8JjTB6cx3X
vh8H25gPF7lqw9hqdXvjGP42xcP0XcYTApMzayluALMjezQTHeHBM2jdShUOjxL2
/tM2v33NoQs6Xx1wKo6w5Bf47R2C8msrwddlqIoznYlaLQbIPfGxs+/yAzEIzczk
IoGtDxRNHl4a1VIqaad48xfOTGbuOVbIooPFqw3+xq8c/EKNaOCaoGvW9qKIT6wD
IOrTV7aSSCXwGJXhfqBby80nV22c5nr1wNsP8xLdoyD5eIEDQBM4LJDmWV4avFpV
wCl4NPdhZlF1j1eLcSSOWXiFxi7SDSO7S6uYMJlIfgawUIrpzQ8/4dmIMNKpbuUQ
3s9121JDgSRO0pwbDtMBgiT/i/ebLwM3P2K/7wjZdfEXzsrTmgTr4zP9BPnp8dp6
cWtwZr+/79iwc38BCQB3cAXOF+03ai3t8BEaOHWDrGqcur1T4QlA4u9f/bg3IYpl
BjnoLm2DNLRc61JS0hP7/w8e/yFsiDpzdYcIowcJMwwidjCVL5waXK1X+R8x32i0
8i+jJr2/TCCkIqIa60uWrB8p0WjMKWTUWDpp5eC4D7FbTJNdFNHq66vIDTph7T/3
0KUZuIlNamluj9/VZxEVMVwdj3sOV24+cjYlyfxC9ARqicyR9wHQKDPcB+Nt8QPS
oaKXQSlhvtk40OtJaGyFK6oBeyNrnOjKEve9rmCl/AxzRjuKdA9jCR3ssUvx2X4q
mun43K6xCiXGxgYD8yt6L2Dl0du/2yD4ZDCc4xRedVlLzJskevA6B1ewPftec3cM
UkbWB70g3ssISUesmh0eI96IsxtuHwtOUzVCIknJan8z2FRU+pAK4REfJnZVWFYy
yUSmwfS8krq0VbB724gTS2xUGI8joiC84+wx+bYmenJLjGpFBDlpmpBNKSaUN/AV
+GuJXgzEamhzChpHmDveIS/puQksT5uehXY8aAR3UdonT6zjZioyKVtDtp7e4g8B
dabg7ZUy8pFYd7ah+8YfKgbysc99zCmKUZAT7iqguM3CwF545sguHRnYQfTjEBk3
uKo0R//pAfMcZsDcaMDHbvpLc8rmo6LWqWt5OsnOh1UTP5nGgSSb6eBCubpeRZ+f
0x2xsUzTNjUEDfnvrAQ+qg==
//pragma protect end_data_block
//pragma protect digest_block
32DvCA7l/2WLhGFmJi5tL83faCM=
//pragma protect end_digest_block
//pragma protect end_protected
