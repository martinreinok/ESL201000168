// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H7YP(K8PDO?D?0)4<EV4-R9MRC<'DGB'%M.FF5G9]"7BB;3W4W"!4SP  
H\[P$/NK1Y6D87=V043"!N@4(XON*X:H_Q@_O8L#FZJZ]4XK6/4EXC   
HPL\ +&HM67(6>.?2/_%WT,#GR_1I9?4A\3R,^M"/7WJZ4MC^(4I@-@  
H[D0L[W!,ZG2/2?JG6FO$"7)M32 =BP\7^&BHEH)/^@MI W/J ;TTR0  
HXXKUKO=4//Z.F)^6N W?'@,H.O4_S4[OS'4=JXFZIY; CZP-781R:P  
`pragma protect encoding=(enctype="uuencode",bytes=6480        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@7QNM29\)QV8$)/M3PKIS[HVS=\EXPQO1+MHR2P)L.(P 
@& 4TWY29#F:?FU???O&T*OA^]&TH,\8( NLS?[_;M?4 
@30"D[L<W7)P4,T/Q54Y7E>5$?2B%.53[AFK6'RJ#B9, 
@!;##:"97GT1TS#1S]^<WVPK F_9,M;):&$SB3+EY1%\ 
@=FV-!J7'A,[Y8QK1XV5XX=8PJ&,1J#$XW&&]8*]R>>@ 
@(LZUXKP70B::X2CL_1CIFX5:C3,'I#$?,OS&_%[38WT 
@GDB@@T)PNLVQDR)YYUS@Y]VX(U8&3P'BJXE]3;S]<%( 
@8B0/_R7@Y\B;,M.VNB>)1\U""YRX#7NA?$\,Y4XP@O0 
@+*6V3D$. 31SN+ Z^@GO=DD12H;2.L3ZD"AT>09Q5@  
@/XXKS. H;]L(.7'V9@9U%VS9>,81,9QZK=0]&D9O <@ 
@*Z;LPZ8(:0\D$X3FMH$\'U2J\(W5T6#9I)^8==;41 X 
@2]55@L)'(M#(4:6N!&8FM,  &A2'KLA##XUJ["H^V;$ 
@B?AZR(3.[0,OJ_G)O^FH$O".(@<Z!0VX#I(3MR0=6UH 
@2IW^ (%&GNG*X58;F KF[+ DVZMVXDRO/.'1*X<);KX 
@*JNVQ?=R+YLEF(/_Y@WB09LTO"-J4_Y$'+?@4>L>;*H 
@R/(!J%4TI7R27S^[/U8!&GP"$.%YLT$:"I8D(9Y=QLP 
@O2+3$\^3B"9793,V?8HICA[E$YBI$X7EAA@\K:8IW9  
@[YXEM22+[DN_3U.$0N/K'5F M*E\N%:VYXD*T:!6[.< 
@3P*4B<(U27N1>;*@ 7?M7,S61Y(5HEHS,MGB=* C:%$ 
@MY*S=G[\[.S0]ME/$<RCD%EVU"G!$"[OO1F)[)]A-(L 
@_R,("9KS7)64PFE[L"AFI5] *V%4 V:]^2\A_;U@5DT 
@OTX542_/NJTD\D?\ZLYZ*EQ^T^DM1ND,I<O-V] 72@P 
@6KB2K;)/6"VZ1V]\Q%H@* AL$.S#CNJ0DE54+9C;.OH 
@$I,4K.Q62A^WO%OL$RRU)(?,84#NI!DADPCF@9)JA'< 
@#7Q4<J'3\DUY[E$%(]:.5=S9>8@]5,M2.?HF\S:P>DX 
@G#ZL2I5-12Z0BR*P(=+2/]?P0!V;[5/#&4]6%5R_EZT 
@B@G\4L>ZA5?>SL;3@]N6*>59'VCI'1Y(L8?M:T6^9Z8 
@>["/DU(VZ=?$+%1L!,W8#$M&4@V.JU<,\=]5;F>/808 
@=-?,XVEC79*"F8 P[\QT6*%Q+L!"K.AMB(3#:ZZ,.:( 
@8#!>#'+QZ8-"W!:,ATSAJ@/L]/GG!.\6<^OJULC_,QD 
@O=7?W7,P'DOAU_6<L+$S$9CM/V751,^G]*D/\M*[1T\ 
@U71$ P+[1L48#GN*LT:@Q4?,4V9@G#LTT\%CE5 5(G$ 
@WUZRO(/UU 9-,X3")V;YO2%/\;HVG%H$JQH47C.'WU( 
@7EH2>P"..K=MDM4@;2?T_928:B8B#XQ\U,0[*A?OOZH 
@>X9*O_I9LX4T 2VB9L9&44;GBK4Z7E@Q$+#UTQ8C-+\ 
@3\IV@ BG>KYS[G^Y6P_LV I+]8E[S\_^G.F"\TNSJ'4 
@!.^61(QANN70/'HO.0.6=DB/;"_T73.ITB18J!#U,&H 
@$'(;3US(HRM4+X>[,0MHKG5^K-SH"0/_1F=6EV?Z=,< 
@1-\HD)!GQR-]@?EZL@RC/-5&@-0D 6!UD;]'ZN=P5L  
@]B=MY:+B?VA6]<;BL%3Y,B;C*L-F$8,?TZ?N"D[[+=4 
@JS!M0V!^&^X*W(+8MO E3[NQV%W;6%H-)1NQ#GK^<6H 
@=ORWBGL0*NA8L2X#:$# ;W) TIUG100[NPC'BFBO6HH 
@O0C":/-BRP=L9Y\CS\W?I0&3]#I5/^+"#*K);IY6T)$ 
@#^:M&F_PU1F&GGBAW 3=K/_]Z'0P,WFV]^"IAF')114 
@X*@?%9E]+@WX2LMAI*3>L')BOD>JTKP,#3@O2898RF@ 
@M+PU'A-K6:^+E I;P7O5OLV]YM3_O8;<>Q@31=)@ZW8 
@NJ>=2FICMN'M92S,B&@Q&F+G5H8\M-+BQ %(L5?*NB@ 
@-+):=2DN'\R'_V<&>F[ AW\:7_93Y"3+LF?Y+G1%6]L 
@VQX? XSAMS.4T!CZ[GA<TT&JJ)9\YQ#YC^F%'(0LU64 
@]O FG4/]\5!)W;5 N%YJ_[M9[!,0;L#X+N3IO; _HJ8 
@<L(58N%'ABO N)[/?9$%X^,4F;;\S=A<-8[U&;V1MT8 
@6'W[DSL&")3.RX XW ?<#(:N?&KVIWM R<[IDLJUX?  
@@&EN)Q@1QA-\@Z+TY6Z&,V*OAGL=[H9H?#2Y7VT.--X 
@Q%,J.*DH*#Y;J7Z7)_@M>I/1(ABM :B-Z9DZJ&OEVJ4 
@U\."=:O&%H$,?#- 5CRTBF%J/V3AM\TJ]N3U.&>_@J$ 
@UDT)0;KUM-]D=UM-5]YO'1_7/9&2]GAYA0(U%&;M^H0 
@_NP.M2::6/: 'QYF-\Z+:5M#\5Q4B*TX!#$K$IGN&), 
@&Y$[0 QJL@_V&(?B0:< N*/8W0M8=B5QSL'K\BT]TSP 
@1FJ&?((3?DJ(I2H(5LHZ0^&P62^4=W4#1XL :Q,X!0X 
@)4SMYDJQ)=<P?U15&VJE:#D2@J:6C/S:MHH7'(304), 
@W@<_;P,WY?P/PP6]SH$N\)H-B:4VY^&XU&/M_'5[AS, 
@]<+#3G:%P_;=+SF3%.0 IR\/7*JY;&K5$]&8+O_VC\L 
@9YDKH:/.0IF=@CM["<5@TRD2)\]!ONEM9O44 &EAG*D 
@N<9Z"M65K7I%Y&(E:1$$$IE3=M<;+@-II+AJV U[QQ< 
@M;!8*_Q@!LCO>QUQH2PD<!8+J9 @FI='F/K$6K]1MT$ 
@CT0]*);F:_>$2^MW.+ DY6=-0FA&(:O06UM0O6!OQS  
@W3S1UKV\7?-X@/T%Z!&G8^J7OV!BFY*L2@HG;KS.E^0 
@AER8.Q4&9:3PS+ETO*D/,SV(9;.(<OZSV)D=S\CXUM, 
@Z4+/!T9<7*MN.TS%4YE>DA7 W,^'\$IB<(=3JK6OPI4 
@*MK)_+_?<O?(B(?VD8K$8*P_Z3P'9E L%EG^8X$+GI( 
@$B3WC2K$W&H$_P;+W,JK2P\08'TZ%Y,G(&*EJ>K2PA< 
@*Q<!HP&>@9;AS,R(=QP01]M8JM,C#)-XN#%#Q\@>TUH 
@*\M [FCTBFT;AEPF]V2]ZP_5Q]FP-Q&T3JKJ!)]:)OX 
@$V> RU"XC%0_/?>@\Z_W]QR[4SM.*Z/^KLZI)M,D[1$ 
@M[F$4J<I7K!=FKS L_P<2XQBIT?-])5?N&1K2NGY/,4 
@C3(]%+6.$^S2(@82ME+VYY8]&IA)5DF^#>^W8%/2[N0 
@0;?K3CKE_&>DKQ_&FN*VWCP-GZZI:W$Q1$!]'+I<.4D 
@!!L7=&AHIHR^0>4O]RV$]U6'%"F_<+J)Y9XWXTYQ.Q@ 
@.?S=,38H4:#R7U'2%++PAD)-JBQA]RV2W)0-(J'^!M$ 
@_Q=\ @^P#* &CFULZRM&'P)?A3W"RCTK;%SY[J6!>JP 
@% S\I=O('8W_?KC'M.U^,6<+C%*#Y.?J2''+UL@B8NX 
@0U+Z%6_#$+?+O-\BM%:?[V)K30TE#9]GC8GY&O02Q:D 
@4$9C+HN.SRE#U7*!H:2JD#RT#VB"?G%&A!;DH4');<P 
@ <=*=OL@TI_N#,G*X%.V_<@L<JS3KG=H>YBD^46CE&( 
@%W GRTBF0K:N:0E@BVZ^]<>KRV5RX%E@(I?:?05^9\\ 
@G-FA?UELZ+$%9:YL(#76I_);I[WT86AG7^KX[N@M 4< 
@2':A=2YZRST 'QF_#9_W7*;]^Z&QA;_[N!B,,@OJ36, 
@D-"$(JZCSD%ATTRWPL9[AYF!Z68V,; 1Q3#HY:R)]-0 
@*NE]_TT(%VWH-2BWX]*#"]Y^M:P&^@XT4]G8>:>V>]P 
@)/; \HL:(9/3H4>4)L=C!*;B?O_GFKFP'FGF#V(EGC@ 
@>G,Z* 9!@,Q8'A;P+V:QV,[7&GOY9L26TR00MZ:E/[0 
@VO%?*]=_=W;MF1Z(Q_1[IDGX46CT,:I<X<80T_H$9:4 
@EB$_/908<;D9@M3+I$LA".Q5Y!;L+<=!I I$8$*:CI( 
@&29Q.0=NIT';&EF>@Q))\6>WX<Y:N)#QE9$KJ;A+<A, 
@"6@EYH&-)K#1(,DEFO_->=&LFT9 0"\WXHEQ[9<&VL\ 
@KH=0B++_=W7U,RL\S^$1.#K.;]G+,<P4B&+\Z=W%XJ@ 
@B&A]P'#"'#PEPEZB5KZ$3[EO>\3N.;7X0:IC!==F-^0 
@_:@C6?+^JXC&77,)>5VY)NT?2CC D(OJ"H2(.>GBVGP 
@>.#Q9FQTYR?ZT)HUWIO9N\W4BH=*,PVT7X#FNGEG8/0 
@A&YC\16D >=<(<>.&L,*PXZ"=(!GS3+\JOK(DH0_:+D 
@<H/76F?]I:QHV9AKJB.-"6IT5#HS4AL&K^#F7DE"=D0 
@U_TOPZTCKE\Q@[.?9UIO\2P4"5L*<29VX7KRWR7D$Q0 
@0<8:!S%8 ZK7[$,"T$$?(+(53!Z:D[MK6[*,EV\__QL 
@H:8&W0)"/OCE1FQL:1?5OOC!N].TR6U](,,;UF,ZJUX 
@UT*C>O;;T="BUG/4"OR<L"KI0&$XHZYGMIM31VH;V*L 
@Q0R&R$Y^G+T*R?0W_/17(8O2=Y#*-KZD]F'!\:!?!8\ 
@ W"Y'U*LR;H#Q.FH;X.SDFJ5UA/(_YF.,=D GK 69L\ 
@@I=]A];GX !DP3<5]S#DOE728CV+*_6BBQG*!%<9]10 
@D=& 0D[H),*WER@)G .\!KHR9G]7-VSYTAY%^\Y8FXH 
@(<TYX]G27?=#Q)0]DYZ26EZ;#CE&TWI816OETM\$O>D 
@/(E=BXU2@\%+>"2NDVU2PS8LLLFG^@6^AB3HU&?2A(< 
@W?MD,EV_P<<(E<*/-69Q! 4O>;"Z/@"6' ]S(9?$23, 
@O13SY8+>JQ]L4K7E_:OS>&'TQEC(^4YT7[>(1_9HY=D 
@GN!!#AT*.7$I</NT@KEOU7&JF.\QEZ8!$*I__9MV+#X 
@LDWR1O4%O?%7Y>^P5N36_^?ZY!5LE.GMRX&^A'D[(], 
@G[6.#SZ?F--A_6S)-<J7#Q_3 86=>W>Y[.:>4#"O#"X 
@VLP#FA]%I]>)1HE*]A05$C-'4[8R_OF94EEB<X15L70 
@?PQZYQIV:F8+^R,;_[4R&"=S81<>:%*9K%+@T;Y,G!< 
@YW_RF")Z+*SG#>^K19PU<Y:-JTS/XP-I[]8+O/^% 78 
@$+S^M;ZCE@R3^=JG_B@$?$WE1+A\D*J5)V\5;%MPCR\ 
@_WLZ+6 4\PE%WW:HBKC39CO?[RLX:5(UF]O++\!.\YL 
@R [[!@[1PJ!\+X>@I61?'=*E& 4&N^4W#( .C:%^?C@ 
@_)Y5Q*?AZ&I903MV 1S,$0[GI/DB_RG7@ /GG7GL=   
@LM5=>VLN:-&L<M:;2#.#R"PP2;;PI#%VQ90!QC8BP>X 
@<SK3DW?VE?(%%Y3T^[.WP=*BB583==)F[^SH:FOUQ3< 
@)O%!RP8H=J/:_UJLLAM?+-P2CZ!/=,]]EX/GJJX!UT, 
@KX/@^5AZ[M.JTT)>6_"XZ#H\J0]$=%O\5N'CL&,C)E< 
@E5!J_7ERDSEGE;H(04-S"(G!?A1R41:9E%$!.)8[J(4 
@+@SK3W/(19$;AO3UJGG%618Z^YKC@'\L]OO^S_GGS], 
@-?,>:HE2X,<M%ZZ&L"6W6:SC/.9[Y4K3VE]./]8!=UP 
@'&[Z\CF?S@\[P @!O8;;JA*M]P073S_SX9^4# ;E&FT 
@]VY\OB"V5.%* ",3P<B9# #I\URZ1I4EY,?]W68XNXP 
@;K1@+ 0Z*$+U1E>[$8ANRL]S5/*T;4XQ7>Q>^0R>,9H 
@0R0<T/J-6\9 %.7]Z- 5\K]<@*>=4,QE!N'CYA8%_5< 
@A\<M#/OS[]:Z-M'?G&;^N+SQOHHWO'&U- C]2)(=T], 
@Y'GCL0#>(6[3T!LO!$('K.LFQ.<M$K8>UEKQKZ-NSX\ 
@JU+5ON)+=?IF"PL1*S+ LV@\@>GA<(-)U\K@/C-T>8, 
@R3)5EXN,H,U:T5H2=TK66O..L-ZBR];#6!RC]Y'Z%&4 
@D,$FT/5_&#\T".ZYTI4/P<7T.'%2Y@(.4SO[4!U/")D 
@_!]FDGTB\PLM2J*4'5_YACH7F#>A_#M18ZB>'L2UK/  
@//8*XGYGPR5,OP-;SACDS*6:&4W.3AB80*U$]W7]%/, 
@0+6?GD8B%JGO*_@,Z?(P3,')IBMD*+HUX'[.F(9()#4 
@/3?P9%[TXGOL2/!S-C0]E]^FSO :N@;38A3#8H]#.:D 
@]7?=N5V6Q=KZU#=JZ4TX5A[!EKF1)SA$&/_&*"Z,;K\ 
@PFL"AZ>)ECGA^!UWP7LC)J>VP9_Y[:7&N'XPI[H$^L@ 
@"=9%QXH!/^"P%F[HU^^5&#A5%E:D;.-I?.)#?>NT@>X 
@L'L>L8RIO_0T2=5B"6T-PI R7?"F&-S4'9USCQ#QED\ 
@9H<,+.Z$D&2Y^<'/'.1,>#GM-D2!56V'][><'#H1^1X 
@.L3Q#>DC!I,Z'I$D+ON?) 3@_$L<DR8\+=+M=%"NN!X 
@@#5<6>F+'L3[;&+*76<SW0J?EQG*(J2'!*) Q:NEIN$ 
@*YFK SVM@^OK;W[*3VU8<07S-TSM%K3(YRK@<@-%"/( 
@7!,TDO.LFR#N#.-BP^2V'8ON.AB>/U2B10-M&7A/PE@ 
@[?]0\QK*^_RU/+EAB5R0J^F#8 ;6S>BSO7LWLN!OB , 
@X3Z.<I0]K1 .N"?<41X][&+R6'BB%Q09B*6JZTVHYG8 
@_"*HU$#'BDG7KZH3U$-FQ%TX%2^J>2?Q=\Y%/,+$_*P 
@=ZCZ57K!:\YNX-ZFU A$M&<]1ZX<[V] G[0P$;-F2A< 
@&FZ\VUDGDOP6LN4"J1-ON1J'5[$\CY^H+[]@C@5$*"4 
@H:R)664QVI=0XBPAX7D67#IZN"'Z7>F[O? &HMV!0:$ 
@!TFBX;P6#)Y9V(F'7"^_1F0V)I.!T"U61\]0>V]C1!T 
@%75_=D#D%^F/_\?BYD7^(@U%*K_BY]A)A4^5UI]@+90 
@:MS[\Y7I/DN/Q7MO?98#V+(T9+0B1"J87MT(;UP)S1< 
@YY;NL;(\G:5+MM:Y0M&QK,V?9&.PI\(S_Q9KL\*GHE4 
@'V4Z?17/Y87)< ?I&'RKK$,"\5S=^F=(Y7!%DU[_[70 
@C$P+]GWDFE/<R?VN]UY#HLYEP%C]2-9CD!DBW%A]_!< 
@@?I,3D3DZ//07SP\*<;Q2Y6E*03KG?^-#0Z,\0Z /ZT 
@&7C@,]=A7(:A4$Q+)!> 6%6LA^36VF$L@R%E$]6P5_\ 
@I=F<_1&(,>U;K64;X"JXDA"[2<OV['.1V9D2^1AY'4@ 
@<-IIE24U+%R&$C%PH16C=,=NL /0>!X1)%XD>OP-=!  
@FI*?>[J-]#O)1+( %"CC4B"O"*M[,VS"9K0OH'9*/+( 
@VK<;(8OLG2Q/RAI)!2 -S'OHA,N,2RH:NF#!8DS&./P 
@LFD@1.F-HSSD7(P59>PXXG/(CI[6VH7M^W1LU_D^I1L 
@DAQ<QHOI"VIR065X*1O70M!V=YN$P(+',0]$@K'G)^X 
@2Z"EMQP?"0T_)9+NQRRYJ/O"[ZSS)W%&##3F1LEM)A\ 
@J3O0: &8#I$*_^W7T'.98TW0!@63)&[R7'+:[5\SV-L 
@4&=V%-#(7<]KU7RQCS"PWWDLFBW1_RGT,U41O7.O-Q8 
@5A0%'570"I69$!4 9^B@]&M[&"]Z*78A+[<Q6\[/V \ 
@.5<NG.&_',8Z9-X?Z"EJ\J5.V&P,=I2AQ-L/Z+O.EWT 
@Q%&JQ8N]-K(\=P"HL4^Z#3+[4D7W:;*P/"P=]:8DEJ4 
@60#DX"+"#/Q?BSG*I]U>1UE0&!95:SX5<W.%H9FS\T$ 
@:D\[$KZKSXI\#06> R6,53O6JU="CJ25>61[S-3@E%X 
@?CG9<-,->X;"0P+G5N#T-H"3&1>T8GJ)@*9<&CI'#J4 
@&=<(5.)&)H_A$BOH]"=!=@3XR@GVLKGZ:=$V([2^.C$ 
@3J4%,AC#QR/T#YCL.N)>&37''N['($FR)@#+B"ARJ%8 
@.E#DH[[2#"!XL!2/^R+']M$T)N)=^/EF89Y\LR"D?I@ 
@N%>78SS9XT$M7)X%M^M-Y;/?0])T1#]>6;*P>H%D*V@ 
@S$%AS/X%U$'@,VUD:E6,O<^/>VE"Z5?IQ3.P:TN@.F0 
@82_^L(E1JX/#@+!)8G\;.D1=I#,);R%*_2>RAX\)++< 
@Q\=I6O:5*SIJZT);)/<\!X0RYS)#ON]GN6^\:MBV[:L 
@+4 4Q.[F!QHE[[ZQ%^?><S_?$?U+4()*21FD]]N9+:\ 
@V\ES#6SC]>K1U5[>+")6#=2>@9'R\.<?6O>+J>:/4!\ 
@KG7*^*!33F82O=0;-Y!YCWQN'>*=$0T7XP:N;J'<,FH 
@!=55'/(S,N.:@?=08+3'T]M5Y=<JR<<@02'C4DC >/P 
@AZ7 E&G1X[TWD9^6+HKQ5;(+F30W&JU4TK M$%X+[5\ 
@JKE*VB-#PG21K]IH<)$I6T=;.7' S:LG2#?EDBUFO[T 
@+S4SE'@5"E=ER60V"RUATGSH AI_.,I4]UQN\4>(O7\ 
@4,?RF-I%((0M YA4(>83S_*\^JK7@;]OG@D'O,::HW( 
@D9R7M8=DBG^<K.LF!2D-6A3RSC+P&K (0.#:^?1#L[( 
@#S184N!LTZSO 5/R\?G( $U#I4,G6T#(_'G7S#@U\,( 
@!VL<#CYGR"YVC096.-5QN-ES,M1Y:G1 :J+X3L8^ !( 
@^O0@O_K3]#8!YBG7;B:?[/R7[PUS[VI,9B^9P&\@0%4 
@;^KDEX"A6;4^B6+5%W1T*B]W@NM7;/)[06\-Y?L59"8 
@3A- =79%7:4$R%Y(=W)YL<7VXW4W?%OC^.F8N4:GS$0 
0<,_F8C/[3R]>RWB1  ;(U@  
`pragma protect end_protected
