// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 03:52:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QVAiwGobQYbVIWy9TKyM4OnqvUPyfkoqiGIAnyHdae0nCRLQojHlUyP5pU11Cj6q
654pnLpstxJIOUXoSBR/8EfgkVzvA1MIEQY5MjUKOpaKWTrsSwAQ/JRG1N78OGmy
U9nF1XZ03Y6wISJ2DGX8Z/ChrStNSEJuSm/PjN/kUSA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13728)
ll1cpHHjU3o9r08r6RcjyycmmAt0ASLIi+qkDUPeoivgWT29wizJuginkE2uypAE
GC14BHfUuHQJ5K55cwFFYd9dOWpF+7/BZ8C4qJsjevgEqQArtciCY5seKsb8cb8E
QzpJz1aENo5mpuD2N1E5pHCYCJJFdI9B8pwLzPMVTEes8tsEwT4dJkG6/UM1cJSX
/BXbegmylzGikV80MyCEhnczb8dsP7DMqzvt0pG5NDBXlhckyDJN4Hn8PI802eWp
qMO9PbzJPoumTQ5yL7xVepTvncgZ6NOUyZFrRmD5QUVfhoqhWrn7us2n48zFO/BL
gWqidDdj2RcdsBK6U+oiwVKZZLkcKYXUF86lDQRQXsNxpiW+wEwCO0uEktnKtPUe
GgnT9U0aU5orLnD1DOl/AqsRnhhmvvdsx49XS4hh253OjzjWk6zwA4vTG/6D4Sgt
v+3CAQ/vs6CofV7TCVzw50D22wuxqt2WePtZF5BkyFBmgDG5/s2W3sQ4Tlb6wH/1
rGT1HdjoBjMKTiANmsvC4IvzxNopiG4plii8mQUIqHN7Keo0DrthGlVzxm6ax2sg
2A6v6+tCtqxYoIcbBUkbnrH/AHy1WDsXRWuRcOxKvtbpDY02SDQE0NxlgHu2sURo
7EHdEx4TyNq+f/C8nJ2Ju+4TyBLTIETrWyNUnQ09mJoSLIMmc8hHLAJRiFFPk5mU
22s0HHqGS9Zx+2N8x6KsqsCyfT0V/4+m/gr8TouV2kuJD0EtWLBETfuSg3FYxSE8
JH4fgA+OEvgDjCyrb2gcRNZ1KfmWKARrTZqs/M12XezxkJ2JuQiMhAQiu+2eckp+
lY44e3p6zx5btt+vhbSCyuqBBePf6Kf2xtZt4eYnMUDnSogkboM/incxNXtKHLsr
1eBc5RXkFlZhgPevIRA7KYpi4TT02OUO/lg/4euRmEtf6RuwCGz50GUhY68H28v5
RZ8PLs4VaiVzmdNHVE/oMJUuxH0KJMthqB0lGriQiycZYueEpyt6rPD6DswztTOU
V7CfXBAblNLVamPt56p/Hlk/xLqPdqJBAyyB9UgAqwDVtu+5zgEJ7nvXIpgDejBN
wGg4L12iiwvNeHCeXgF4/EAmbde+0Anh1vNzvKcvRJt5P3EOwMrDbymBi7MGqEFl
/MMvQgouXUeOAplrg3HGXKsD9QU130Urkl2hy0YGhLBCXEroDNn9MpVyM4AveiDF
ttsd8Ne8f5yYtXCMq/VR/5M/6eKZMCrmwtsACCVlV8QOUJuSxa5f+LGSEXdTdotj
+ZpYJA4c0LE3sPRMaAH9J1xgpvAZhzybkwYveJ2L05JHYFxH4f0WbodVg3qfZGiY
u8sSh6munEFCA1noO/ayr64FggcHmorDD9p5sBbMuDsMc31058X0lQcbTAeMFcnP
hkWHs5+WMXT93iPub4WD5beHsiepWgUPEHqHFZkY0lf4vAPuIAVIWruC3CNLRTze
rbe0Ihg3panXo/vInPjDL9hwHV889luQ3D4Zf67Qhpx1WZZAgdI111UvN+tNcoSy
rs9YPt3aqhfnkwDFrcElMoo5zWF7YqNgn0+VJZdgLWGACBHaXoTN7QSTZaB8CkqM
QXiw275JZP87uW4kYkHcIMw6dL9Sv6GNTkFttsltbgFIrunUaKOB7iuwmz1HuMVa
3fo5E9yiTzNbtDhGkUZpVBMjFXZb/E9sMdWzpLce+WLEiqpTeYMgeq6GUrGSSH0Z
TDvZLeQW7ZB+7qV+N8GX6ohMSuqnfwbxv/ixKbsHhzky87BnReOYi4Mk4RfUHduO
IMlbY4Af1qEoWgPnFwQn9mLCiatcF5IFX6g8UeqZ9cQ7lMXdWkJKqKrXd+hc0A1+
fU9Tmbkpkhk9wGTrZV9WDYqZBPlEfFfzQsnOZIluTQc1H1v1Abpac3fZOu+y8DPI
bsggE5edXJBlkr7qftUPJlfoFU5nwqHo9xhsDM4UjJLfm4U9wI/LwBJKq0TnpRRg
02/OhDIGn0Sm9w6ks+NOnSgrlWyRzv1u4b6SAcm3vUWH4fkjZRFVJnev2MZyL572
EV7pIs3yS34E1aY1S6XYz/d+kRmeqlfcm2n1urpPlZuJGdhEiL3I5TaC8T1YkGFi
7k8hoAvnPQZxL+02FUGNdtLCqL9r+iRIYZ5YJQdRBWTVWvtCAYvHZeYkPy1aQstv
cCXTf5ZKWJb7Nh+kM/8Tu9Qyqzj3/fQn4q7bWKpkZ8aJNHebJguupSrcYZDMiT1i
kN1w0W35ylM4z+mbBvY3dGwf87QNTh2U63/DqLpF8xATEmgSUJuyJr7ZtURf/ZwU
lXJrb7pU5DayMvYd2NWKuMwMdVXOF8LmP4TpobC6vfX36Zx3K4kRlTqiVgwfCFQd
dWjQ1a//dTVZJs6Xg3p9Em9xnMd2cfEHFoyUgh5y7NdGDfShxOWipS71eoih6cvg
ImicIh4ipuBmO3OFYnJ874uu76IWCAFI1TVDNmBwysxKMAlxpLuENQjd1XlefV+s
mCMJRGAqxvV4P4ChnsQE9Q0CTsCy4RSZE15mGYIBS0ZEZusEsIXCvW7hZoFs5MWX
JlHLRtO28qmqcJPGD4bjpgIpG1iLarQIcdYPVTpg1P3vrlW/aK+LNQeLz2oHTO5M
LVDB/bhiDA9Cyo+QscSbuKt0kKpAXUnXnV4VXPaiDYNet+f2SQ+im4pLAI94cISn
VW2LM2BYbMpfUlLHf1FGLsUAqTqBLmwuOM2fYFzJSMo9O3PVEV/8uoCW6Uhl6bEM
Q/arxHrL3IDCOWasdBDyKxvQf0n/MHgpSiBSaooJFLwAjd92kE9wjoCx89GNd0aV
shMel83bXbVGk8u9v+FCpoUH4TfRPBHttuJIEhUVQ5sNylRjApRiDtCA9UYsze+X
Jr7n5YC00BGoJy1zHnG8FbKkDpdsMwHtVmPvbu6I3rMhSKJEDNhayhlOvojysAps
PFpppUSnf5AioQYyu5xx8iooqjFkCv63604a7rUoiYPJdQJ1Dtp2izy5SM9Tq73o
C2Vp9g6ZDTRfJYURNeVskI6tDv1eTmFxTTIJeN6/F3X07RmsBp1BZoK+qlsAvHK5
OyqomZ7LAQQBAYGI1yrMhhxCiCUvJ6bXPhssDdgvth2HCNdh3KkQQaTrVeoPODcS
ql5wZVHzuGXVoSBTxLx/APvHM4i10bhQWMOx1KcaHjrfcuaTf1Nj+IwzfcgKDrN8
Ec0qxNHZZ++qsjAkZCYzdnS17VEVqrw65zNmrlptXMtYRn/kglk7wuVj8uhwTuqf
/cp8qp/YRYgg2tHDfgbAe18mDBxBUf9ZQTWmuSjeOVBxHXNTLDX5RnjuYAWNQCP4
7Dyld+6Dsz8heTWyZodt9ntg3vVosbWS4AVZUa4Z2jHd5/wnpgnX8XZKiWak9pKl
kYiIS/qpTYNtY5bTnlm88tEDvITH2KEa6wb0ZcPNupNzEy5gM2Ywqm8BiG8y31rS
Evl0AVmsd5OHoBDQ6hS98QDI7AYafE6/QzMQvkKLTrTgPz0ADmXSEiopUTD4JmmX
Qp26hNVFyIHW1J6mycbpl3kmEDw79rlZXYjOq+kMUMvGjKVRpD8RLC7NyLMABeZS
U5I/rSBBduAzIvGzDIFG3FZCvQm1Yd9yIap7M4K1LFnTrf1ctSM4+FS2ye6uIAwA
R21AAC23HxUZGQaUdxq/PIvMpynhLCGgkMNdHk59R8hxXknUn3SQAdvDjcrYdbsH
rC8UQI4yj4iOumNO8LK9jOR6gW2G1HJzy+MB6DqIrzjQ8pmLOU69zKEXWNvs07FM
Fz3d6KU57pqGxP9Fel9aFTpKB/vru6f5qrt4Y+yKa4wKMGMuXVVMsMGiNthf0Agz
BaYCfRr0bchQRVqBcItV09xJ0eET9v+Xw3V38lHX2auKN0vTYC2wceeTZq1r5H4Y
TIu3F+lmxGlq+SiLXvuOQr100SnIoP2k8oYGwRiizA7LawN8dQepJ7SqkUTbY2On
nrv6fUtEYHx5JtRWxuvje1yyTEeLWC29QFmTeaLgyHBhAMZ5QehD5lf1AiF5OUDt
z8CH9k90jmbD6NYHGB7PrudtlETo9oReHWEnypT6H5Tz0j5RcwN8UukA6ZFQh/LN
zIoNI35fVLikDIp+0ZM9tkCH/2JKKhDzBFyyeyic8bow636W3wV5Gws3lXgbCzsb
wZAPTIlnZUUcpt2+wloo4XbU4xLOrobyRY8EF21R6c9SpkI5EHkHEJO6sAuWQleP
5HnIuMMAF8xGhhXTbSRLObtasECw7Oxo3voI+INr/9K092CMIMD5KYNpIrdvbDzh
tmrAUoJL1ghxKG1avvN4mhqEejAT5RGqe74TYgIPifduw5DVGNTgcLiWsypGe+hY
Tl+yTSNYHYFukFk+wAe6P42mtZfrav6tpwa73b8OyKDHXa7EOzihg41Y7hgmZrO8
aowqMmwFE/6XvQ+BLBc0Gncbpn4WzpO6jS4m/GSe1suoS6hB5MKOjlTJ8xIPjzw4
+0L6vx8wdlDZ1copA2wLZ3FMjkuD1ew2AjIJjNvtdz4Bcig+5YqIFZd80ht0mRoR
DsY3il7qhTxes4p/oxn7gkeUwhkFR31IQXDPeBvAJQKJf4KIyk+6TfM46Wu7GnIT
CB0d4T3mgbDknZkWISchSHqsNup/RkNgAzfDwn4ZoplWNPZStQlpl9MOrjLNFAJ2
A9lF4HLNr8UT1Lqfo5u1mk5CbXVryIJL5h7RwQWEk7yY+BM+Rhe9XrXNUtvnmOIj
cF0J8/MdACc0x6JypOYtDu2MNP5GMRKCzhW4S4K/sleecRCBPMitWrt9lnry2iEP
Obgc4Sr/urwm2MyJLsA4mP9Ri+F3ZwEQYeR+gcl6CP9vFH+5KLPlI0oNZi89SVlN
sVeM9rQqdh/Z+V2lIcHHALUrdTnBJg9DTznBtJ72nBDvUsO631fyHwsdy1RM5ct4
Z/6AYTcODlUhn9F/x/bAk5K1WOwh2C1uvZwPPa40Ok14JHBosfTst5Eb6RIZl6o6
SD00WDxH68JVfldw3EuHgWzyhSs3F3YkG8yl2dN4tYuwNrce3VCshtLifvhjtC/0
HNW4ZabNDVTIm3lxy7Pvs3BkmqTVue1BZJk4sOvXNNa5LhmvwlUovDCcqXwfkD7r
JKp851ghH+i3Lm82Xg4Iu7pLARWcn5u0yDCp3F4X84iBzAO3E+oAU7lQTeFwWGaS
YKd9W4ZT18aimuhyrb5AdrYerJ11pAXG4oGRjJ6wEK1Syq0vBJ6iqn6k86nIjzeA
MTMip+6yNutDkFw01lwABE4/BYkqDgZ6tUGiNIAbSvmR2IwiyNaoGJU0rtO8Onp/
b9ICZYX52rbyA1tLhiolgkz2bF8Gd9dUqd3LpdgFjYpEmgQzoR4M0A/yya+Y27DO
pGqc76mPNhyvN9uB/OsEl32AjOuIHtbcG2oC7DUY4UaiblJ/xkRWTKmpS8nseyUD
rpQkSdRA8ZwlAAl/l150W85aAvrDMI//7hAyfwrAQY3IEDC8f7t7l65jAZ4YsXEY
7YDcmK33tkmTRMJgq4q1/7xHeZgYDazQpIhuDmKfGsP/GxlvX0QNDZJjEyJpdTyZ
cMfUzdgLK/5IfOPF/BE+XkUgv+ZJgU44oxE1X0NdnM93Wvza4TUT2wVesTXbkYQa
XX5Sew4Y1uJZ/UvcCs4z+74WmoZrqtXy18a8rBpyVJCRBao3uOvsemQpyNk/Y2WN
BZ4+5atCW+8iIP2N1GDJczT4Qni2kW6Spq8LfXmUp6kuWBAnVzXameTIsMbgp6ln
v5i0J0JP2UTX2msFG48l1wpmC6BQlIxf/FT0Kthi2BspX9DxvIG1nXQgYHN9oHou
STe1dIZQEEV1KzCrLFsDMiywPfs9TsyJITpJ02diNryp6edM3ZpUSO7cE2b9KBhb
LdkwLh6wt2qCyLV7iZ6IJSgsauUyx1teVnPlY0/aqQ4Dc/xUIqVkWqFuTAUr9T3L
Gvv1JoaEZqoaO/bT+dUoejDLmhtse5tWwjTNpb310g6HObcgQANaY2fbYnWIP7ih
0LsqurfveWnSqj7pIPiIuT1ttVt54JrTNrbHKIjUyQxKthuNClR+jeiOzy8rmelD
ntNqMdMHYUpTzlBZ95h0YS+LOx51dxF+0yO2bzlC+Q1wA7o3yfiNL89j7KlCRzvi
6KsPtyYsSO8Dpa00VCVJmqgAs3lMhkglbEHOc4vmMQQND/mHcPe9itCT30cJHkbd
BmPigACcCYDC5tEay7nKDIkuV1ni2Jv1FOrvw3N65OGNPq4gHe009pv2NOJYT3zt
qJHni5jEPoBPIkXxqh3knELVNLu/tL92etQ0CC6wfgXEH2aCqDHITA+XhPpeJY5/
bjCJ9rXWQaDuSO4P7XBo6OLkRC5ZLTulkJd3zimvIW41Gi1COxFqurcJlwKG/RUg
AEUrC/KUSm5m/iRLO2mc9LvQgT8l6dpDAHdsWdBx2UY7fXCVAXjtAzncexPKboQ0
P2H0Ed7HpPjl4SuIqJqtiTRRQjcZMFLoVDRcm1JdnZ4Za4IgLa4HtGt41PGS1Hfu
lQd7nxR7JcTzFthw6PUtc4zyzet+BArQEOQZ7rqWIgwMAUOGfBFgGG589Z7/XSb0
3euOnHcO+r3qDJJGtG+yKyLfp6X5R/eHAIgD+Ovxj0b8/00qcNj/HJI/tMjVjuSW
/9vjNmkuQhQvR//VnErwzTxnC9jRHOebkvjKMntCJpFcoaOqAAx6C/5wthJroUEJ
CP4RvpHrySWeDkjLxBG8cJWdOOpwXIwnaTqmKVxoJFPzubdZ1T4CWBzUivTtvRfZ
YvNGjlJfc9ndvTkd7c06xDFEjtaZ2c1F7MCe2uGFByh86b6YLWqKHgf00n57mq3x
0hg/HYNHvsQYGmyrnNQpdq9Znh8vnOKKDZuuh2Vlro4PGBpvIpoTInrBhn3NaKpE
tYXgSOb3iT52VuAaGzebPKhSGUhXjTNHSHxP/HTzzHdgwjJUJkzgVp//APHM3s6K
ZnFqvdJb4fK8eobTkLTm/DXX5oX6U6Lf/ShMcdQ1WvGPuO8JCXkpAqBzKE2NBpUL
P1woBr9U62MuFGZUrzurjBg8cRVHDBmbZ/X4ZFS9zUCAhxCaakptfuYLP+P/WYW0
zbZ7V/hYrVGsnBz94UCBmGWi08lhwvmechsvj2KPtxDWLvcN+lroNzuPl0dafRT4
oJiB8vMAEFDkxRMkz1wrV8aoCek9TtrTzWCQ5slya14AV91M05l72hYPEaDuyBls
uD6+kqda5ZYswtk+Yf75Jz7fAKCn+aYb8kdcX+tLDv7rjGHygaAet/2Sf6ZttIid
Z2OayAtKlBq66IL6o1jAooCettsw2Kvp+/YqJ22PxgB1LxJzjPAIsr142rbOZ5vk
7MHsYqvdgP5ifrxi5s8n4efZ/3AJPviGVhOasMf5L4Id8JbdQm4dDp+tX+yUgsIL
SEnVSmelCE79lRE3l3xdPZlPhsyF9VK+Hsx/YSSVatUxEwlRDPYICL0AK1QuMeJK
34OSGTYdRHKrVou8FHq50Ke4O3MHLVkRSa/hKakdzpLDAM39W0pF3Mk8Hu+ZWNsy
gHdFrdsB1wcxnQtCCtBvqmEKgfkcOprLJDJ3EZTGqHQU8HNcuwxjDMDgSgdkbPy/
yAvJzzGMYLz4y+bVcPcrKvYVJYxhj2oA+UCJY/NDCrnJ6/XxzrMTu/suvoXcRYWk
qqoEtZwMCZKc/ft8QYppMB4k+rg8dKInvCJEvrkNnpC4wvP3QfNoxBGBnoJ3uQng
qFCjYOdy36aaN85ecyx28wrCPGYYEw/drssQp3LCfdyzCj5pWYknC5bHLk6q9fHt
gft+3teq+ZamBi9rr7EclyxESAWlMVcR2bQkyRa9vcgChGkeirwvpnkyEdlD9X3y
OlSSexScXSan6Da7T2ozr7TlTWJSED7KQfatjP5GyoWgzCrPc4l7x+Rc59XR5Mj9
VxWEwPpacLrbjpOb1xp/7DwaH3ucqkwcv5kNb2ALrZEVSQ9/nLSpYrJyvqTP04Go
Y769ILmFt6UgCUMSj7EzTJgrV/lFhEGm+M2EkDgEpBVRvrytNMvJJYDR73r9xZhM
1SI8nEsDinDAGY7xvIQ012BEI59+77mJqR4vu31Xz4g4rGCaJ4npUqR26qHeiR1H
kgCJB5ZeG1GvsZjQSR1vmKm3V4gPdJBLfyReufskwr2nmbutb0/s2jyZxgGmGPFJ
Vc4SPFdR8XZCYeMtUPDTYo/dORFSjU/NnTz/St05XFVXC4XntioCkjz3iGZTZRkG
Q4DTvACFN+1rj1hU4pTjxwZj2GlgCDmEOmlk/FYxbZ0aFsGomWiIMmM3J4xBCMru
8lL89kVGZDEKFxl1gwEKXiro4x4BCdl+QZOQ8WTFFZQL/pdB+ZPcHxbcGyefqsTi
gQ983dPiL9AtZDVOU0mGl35xBJGK/NQRF3PtUOLASZua77jbvOH6rF0f7+Myk345
7ZKWrwX3BP1hkzEkrYSarg+NJqhjWqv+aiH9BvHIZIsJO9dAJnGoS4PJmBQEtlwP
bqOJfRpuSdiB8elmOlfC3+GdH7JY4KY+djUbtcmENF3bPY/0QH1Uc1rNZYFB9IBW
P//jCkwvGHFoFOj8L7fWvXPXZMLhiMXvanNH/bm6zrJ6yGvmD+T66D0iXZrEwpdV
kixy/64oTptagI03ns7zou0EpwocEhZoizGPhYyxmg3+/bzcKYlj5b6+b5AFSD7f
r3riJHStWG9uKzh/b4+ZLnSTCWDGysOobum9lA0kU579UYjbRAaTSWhYyzXD487/
MSy63132opUiPaD1w07JUvZXIrfGMLCHJpqCAmtAMcEw2Yy9yOOml1926nYmzuNV
aOV2pxIApNxa151AJwK9aaOPpy3ZGvwXME1jTjSZIMHJA2GUafqv4qV/1g2TX0S9
HxUy0VhRyDo9ZWAn1TRe7OTSNLXj7iGcO887p8vtI+KZwxiLoRmaf/quUGW9fFqy
P9hTHQv3apgww8lAadOje3JnioJ7ICquVL9jA7NUmWy+wlOw4413IRkTczXj7E4M
jMiRifAVFXY2pzb74mhZCFzLenYGWisbzAs7/IjTVNq5l+PU06wGRI+Z2zzenaQv
GrSAOMX4KtHpCTP5WDStzFGero0sKRlPV7FGnmzMJTCH6QiyUIxMrfmUAFmVehqS
4TlgXXKoTVybH8bloZJbnmQtbtwwZO0ChaJ0PPlOwWlWUSgT+bSbmqzdeMdMsGKX
ezyYM2kPyN09GIPxSj8wSVLshQZ6upov4O+Ik1sQ2PZ0oaMQkD4sd4wXmpZx3HFd
CBrz/0SfAK+0+T9HBzDvTVR2TyJxjRpfSbN+oOq1bmpckDSbeeGpu/zgXdUPMW0A
NZXuUgmZKw+pNMVSAtc1DsVkk1B9tY5ZwRNjc2k93H3tCNqoXAD/vzpNakNH8WCY
ioZuxGvkJwvmedgMm+JKxHoYkVXq5IbvREUgniZOxNtTbMd42QaA1O9N1LBLCa3S
zUIAs3n9Dxxw8kNSl6Fzb4y+AWR0jaURRa9MQxOKmwUeYa/NKchZPbE3ZqLp3K48
p6j9vYlTqBNyfZYSqg1Yke0mcOrrlTesTIPmH47bMuZyUlUVfFRKzQJ14oRVwf7I
HKImhlT/DF/c4G8evRaG0608PP549OdUkM8y13UhUGwP/nNIUlap2jtV2PRfaSNd
iBwTvSo+yYYTbMs6TQ5NFloEYkF904rQzmb9N6evpW3B2D19Wg1rgKQvK9OilSpg
lLDhym49Ojn8foZdvD03TTC4/RykGQ0NZzhg2tBak3L6yh+HrCVa56t+MF06A/Ax
XLERfpimpmzr61LAQubeSSQ915DrSteONwPHfqKlLYc6gSwOdvxKVjLl9nsudVXT
zIo7q7Z2Ghcti2v7rFUlp3VEGSj/m9ajh80Vks8iLO/itcEJ+IThP8ZRFpwkyY+G
D8LPgqh533b1N76cmqaG483j86pYuQpRb9yey9RDn21LfjmZYqdFxeXzNHWbS2mb
xLdh6V73owAPDjLLWfhuM+RZnzjNs5l2gWNDcTZuK5MtGx5b5Qmw0Cqaa19CvssY
wMP6Q3mWMjFSrdRK1PuR2qoy+DNTB/jVIXniR6B5ollfzOXefwQfzpVDMc0WNswx
avMbG+d8Bnc3S6oCUO5pf3pSixhKRl/2cy6rdKuSOnoDx2sVRC6yn/LUIjagXn6P
zSyyK3Zw+VaJNtE3IsYVBbo8eg950KFbVB2CtDaQ5+sheN50TtSh91dCsD7YOkd1
MX/lyk/ppYS8ofGXh+Z+SziAAymMpcDxITfO8m523FtrdkGGx2CIQs/tLm/s64zu
2QZ/uHesnNu0ZyUmd4tm+qO9PuNzb0ur6tA4zaCIBqHPOwzluIn8rPnlLkAJ9sai
UU5sKHe6kHKdYEMy5riK3tcKrBNE6Tbjz5EKp4nSqermM6zOQDsYYPCf3sdQQo1t
4PuUCoCST4iTwneVQUfQyKN5vsnQHZaLIjbhiv14Dzp7xdXwBoY2veNiniwHniBa
i32gwNRHuZk1rbRQMVfInuhvMHt6kN9POzyRBjqJVcAWkidHzJG8bE1C5VOHIn4l
xmWkjgjkI5Dzx55yMd9TWV2oNWhTutHIsjXZZ5yk6a3o9JAYiG1SeO9myW1jsZb0
hKCt9ij5MvpUXeo0RuZkmdALigVmxtR+yzxJktzlyIPs5kymwLJ1aGRWzeV7ARvR
Wi7VwC+VMFvdioe/KLAbPFg7qUpYgiMo8TTC1iDSLZBMVc/1vThO5rZOKEK94pRh
yvLuccZr80N2sTlYjOUBLPWP2h1YHGZoXk7mxidGTHeH1TjkyDjvpse+k8SP3DxD
8sB5QjcrlgW1mj2SlQ8QwZynrg8rTWErPQqexN6eHHerdJsLV81TvBtwcF5CIpuC
ni7n6x8/YWgJJSqnKD8vIqlQW5ggfmuRxIkWr/FqbyFRAncR9Oqy66ofURBCbpmE
Qqp2Y08ulxQKW9/EOebfjmYoqjZf7AHS1s5lyshvydSj4Afv4CO1B5QybE1nlKIU
Xu92bAZ9h6kn10WxR0JmBjlxDW2hv1AGPdFVZWE3gy1DxlJfnWCCrp27Szu8thHE
Z5XY0q/TUaNtCY4oIEmBmi+b+k5xfGlGtjJxOrwO8mZ7ZrdAeF9W+D3qSux18Pl4
Sqgo1q+/VpPwiG1FaLzbQrhRCjUH7aY3JfaiLhs2oMrZU5Q1S7PAwgDwUpL/5Klj
BYXvxN2XYaH+brPOdcSVwFKy9IEei3JhFuqcVugVDOY+gGIFDox1w1b+IsYlDWbv
p/AQ2buWQ4GWxIPSWyBXtgr9bx9LcyRkeL2Kg0o14G7eniIfKXYnXAY8i6ArlyMm
gIw2ayWpf5ZrAdOZLQdY/+Csr5Veva3Q6mEoj1QfNhu3+okMLvFqnnIEex0x5GOg
uwQzNvhl4r3bCdlC3TBCx8EL3mXcy2FRj1ZIV6LNtdHgb6GLV/j4BupungCNBP7Z
qI++E5I5IPVJVkM8dskYqq5i3l+99xpCAc/64iFHxq8zWEVpDUNqrgPNT/CbyBeN
rfTAGO9qrCKfliGECQmEeOUb2YZbyNqD4n8s2OHLOHwPI3l1HpBrs+RRMQP/GUEb
xkY9zmqwx/QqwgblcTx0gU7+biJEdl+hRcJwKgeywFHC5s2OzSTP28Kypn4TqviK
CjNYc0uQLsOJFJaJfOyihE2PHTU1OI7CqmQss67ZCL5dWnnD1pOkfy3xY0S+309g
JKxG2Niz54V4uybUjoU3WdDAnx+HNNJLfByI0UwqNsZ8wj2yAkb7BS6G3GcEEF6O
HhIgaS4Yu4SYxfBvU2LUy8coi+8RxY3wMRG23gmQnG7Z5fxrceQclnzN80k/pgvh
Y4GeFa3ymLLdcA3ezoPoLP7cKh+ajaeQ/qeJphPhyhQNgELCdzmQG5kQ8UBbTFEX
bPyuegdJDfYpuuRUJngiizLYKVtlGtdeTieb3RhRYbm5ySw7TAIDWon3mPqV40mH
w4+BGqpXpcQFKrUbUW7gvVVoP9v5A5HPzUshwjmGR+J3xtmq58DldLmrob7XHfq5
MovynSObJdzk9n61opjgmwxJfCiKE9Sy9Bfnw/3SBSIzo3FyFVRm8ZdliBojRw9X
ofovIq85vfziVrWtZFOV08FR0/YCl++PlTLis1O5wiuFm4cEhMNHQYdZgv0oLKu2
28Uji9eLAX49tXbAhmz98OPsTFC3fccJTrBtVw1aNCHO3n4od1exKk6PVrceqJ37
7of1Mhq+zYSZOLMTOeVGgrIHnQfRZA+rkcccEMiICXM0cX6/6vk3KrbfTQu/P8yV
w6pBRnmt4KhMIX6cfQsTgGcSmT8g1MkUDL8vJHLW4LVEh+FdirTPVG7btarC+8cI
nTaP7HlZqCYyhjSW4RI6wqw2XBQPyzFLv3oWdBlyjoMlp8jVJZt/d7D3pWWW5FrY
Pk98xkBHIeSEXQU5FaqEfACouLFKZX1Pm6LCbcYT+kwoweUDighoLzU8TcKCuZzV
rTDtYLOEPAtP3KibzRPvtnLiz4jLcpa4PeRUaYGquJSc5nwH8QjeJ4E/f+1uuEvj
lIr7PUD+CP7h0bLreBPELX/LW9r1j9yrbCesRRbKkGQmdFwpDzyWUuPupp3SKkU9
FlG+ZSHQtribEdWhQhFgIiANZ18LMnuTnksuYFFtyM9uu4cydFznwjMiSc+aeFhf
9aYFBFBE/8VOkdSBdy75K57LVTJdvoT0ltJXMQsYsoaSONpyw68JZfHfFIwRpyCt
fw5VHkhms6AW+s6pC7ifMw6gFbzqzV8usix5HSgZBO24K2Qr8e6HGIUKaWHXLdIP
SubEUQpWCxJxtc5rdjbJGnnlBa4vqJt7AmiWVE9z+mzoRDgtpwswl5El+xbNtR3B
HTtoR6ZXkE/NPwcoU+r5CwRXPERlLCTzuWJh6MtC2oRQ54G6lkCbMtGkhrQSXqFo
CHLGERdvkGcNVGv1eusSGGufPjyC7BHTsZ9CV5apDMTUp87e8KewXwA1cf/RN7Gu
e+lqrktQds7Yn+c9z/EWd7c4Yh+p8iP4K/E4FpoCK8rpuxhAVevrpnyH069i+oPY
99eioyUMB8R6ICesn4HRf2Vs7HBmsXeDNf0ZwX+SAD9phbxGUBUgprNu81vZ7y8J
edGHpf0gQx2ebauGsufPDmAhOThRGE2aDsBBHAH/QIQonNOy+J+ePVaqCLL1uf8L
Z/mRaWP+Lpn7nWmpmKYTdhsFOwnxQAWHPSq49yeaPD/GpK5j4brjQXrn1X+azy4M
anu/RqapjlRL9ceUfXuMYQtak3ECkgugDqvQrvhe7DymRTHmI2MbkeR32jx2p2MA
3J7HMskP2Q+1nMWl+mI9pexn222GFcmQe7Xc7Ct+gYHINR94AZ4nUstbrjidv9Qe
XjK1/UycXbZIEGAvYDd3OfyhziFvd19EZMdqPs3rJfx5pKlxDp5/2odP2zz29wQz
7d2j9YV6kBqmcjiaC7DSCHz7jNVJIUdegLO5CT4y3Lt/3BdepNmvPRlTlyImp89f
U6rLC9KtwfnSvdSM4L03jLKz60+6nVulyIJuhSJw/7sPx8ov95kBozd6XHO7l9XJ
viPMS56P0PWivtvGt+auXdPAg3+tXxW1W+rjb1jY+0I6dOytGJrJgcXHBCezZrrv
j97zyQWkBj1piAjBFwHEqIeqvMxWtWxHY1FAcD8V82qaYYXeOhXRNLik1tO9yBG+
dSWOKE9ktovDWWK9buvfRo5VlttkSX2UvjiAIaRWXhraW6/yIw2zaX3UcPusRzoe
YAy1CUXHV7Pbp+wYQlxUt5wVjoI9mVt142mfS9QAYci4GCSKvY58HQWNPFQndg9Q
XKQFpF3rXu0E/LX/SFbO/2ASVS0DZ2wMccdOEhLplnan5t5IUc0vgtivvBV2X72i
HXXwu8rKnXVo0pkq0a1UhG+yx3S9CAYS5Y5dXJ6qHGNKPdnX7nNHFl3W3H/e/otr
qSqyeU7S0Uq62AVLAeCBpS6G1Eig6rI/Mi6zH/bmr1EZLcpZJwOoiYtOTdamq4by
mscUeE1c9T/5Y7BMZhsAacoFOD0YnYuXdc0BSRlnCpcEL1pdhTg67qo6KoRIx+uA
jo8JYYG0RMUheOKVIYK/L4oY5qXKyZnwM9vkkCyrixBtsSb/G3nLKobEsm6vnXzQ
nfPBOsOKEza4mVhC9puCIaLAV69ZpZhHj7/RLyU1Zc/VJELwdGCBzkRmU+LG6VO2
kPLCWd8h0MK+DiRVXbylqLHFEFWkesSQSm7cOY0jqPkBfqp46ZjArtEVXLbI+/rc
PQKkWiO1DSoOP327Bfo0b4rYZcXbLzFsRXAHcncX2Fw20B3KLZMlHkCgEVRZsGw7
H3yZqEVqgr1rdM7qaElVvhK1xNyUDWNWo6V5hgpAHJaBos1HlhGVdsBxot32ae56
JUpWxhR/iuF0E+Sx53SXUChjgrRA5BVy1+EPU+wHvsQfMjGFTTG3xWDkKSrnijdq
2fg+btYwHUVgBJlPXZy1I5jycnYdYRQKDBZaaUlGtUUdYP1u9VyQYsfU3ZvEoF+p
Wd6BYUcR1l03nrg/ee/MszI0SMQvAcb3xLUYmH/Ux4WB5iq67CNrCpaLE4z+pKTz
VaxnnOEWWUiDmWmba5rGRSve8znn1hxz0X4odV0sZhub4EDNgt8kwyFxP/mPKjCt
Ht7PibfVwrK9WjrIXgo7hFOLXdJFsOs9HRrrA+kF0tZCqjScc/7cJnQgEvlrdzME
1uRvqC/GVVlpvmhzZ7y5GVEhgrBZqduMxr/Q495La8OPXBZmMwZ/Bl0ISvBtXpdK
AT5H0GAv45nii2EnDkPfyEDS22/XRuWeeCVRJY128tdAqgVe2qQAJHLbaExdod7h
k+Dch5ZYAvixdCrhsi5T2pCiCIbQyXAyT+ucPeH/QY8W2estt42xOAZoMISMlFP8
eu5hLQqz/dhsOpw7V07uPb1DwUlVX3/zsiAEp2ZZ6QRI+5jASHeNCeQezKnizR8c
FxnXQbtIm621ygjAFUBMFqPf/91JdiWewFVOE6cOWWgLDw4pZwGBHXwbKsANCbB/
dPNjAxIsRfwmNst2X+OU9F4p2Iw8PIFNXm+OtecWA9Tieb/UVKxesNbUCIQikl1z
dSMfSbrV/c7CPnoPBAgqE2SLX8i3MUpr8ULlMXuexVurUJV8aGuemv34LQHLn24A
MwZ0fmlGU6OqnKgGXMPoN4nnNr3lBTlgteHE9Pqnl7WJYjymMPAvP4llSIwI+0Hl
39EButMzs+CZ7PyavHUrABFLji8qcNkibiubqAAwt3KDNyeLV2E4KJP8YmRPXJak
/oWFZr4W5ITtj/r3tkXliJeScgyD0XVEM2fOesOYvTc1F3oQBFjKv3ezFN427IJS
ib+FrQyL6OrI2HSRvy08dYbYEh9UfQGRHHQMO1p2BBCr2A2Z3l8oKqpLb4BV6TPH
iOuDSr82428JM0emv8Jdp3pIQqzEdG9pWUMAECQYFxiXNjrNoXukL/BqL/MMZmLy
ct7XNrHtCsh2GEaIr+i+UkZfySvj8XLRDiz8Rlha+UAzLVDa2LL77Sm36tpf6jPc
WOlHk7018KurQ3PA3bp568Fz5oj8dLkDdypQTE1KNETpflwyg3rZHDLk9DYMMWEB
md1YXsY4la9v7cC6dG3geEQdpbfh38Y5LexzTEDvU8DGDutKgSA/41p7x9pH1LiZ
6ph/9UUUDeVLyyHbjTooLmYAa2+G7TF+Z718UsN9MEfhoI0fGQBclYCuZ0PcOqiQ
dtaqSczK2/41e+RbiU6R+LQ2TqrEXzHl2UWZB4VoLhRUGR8OyJGW3j0mOPRDISKI
RBXOIJtjNc8pkI0focppANjZxR/Ij6XOspptM5zjodYBKX/1nquqGP9bodxoZjfg
Zj2ZgjjUlR6aTlj1YUxSe66ejjGWkPCnH0dWUDqrVCh+c1FPGI/Nd2GqZqi7FIcs
gI8VTvrGfqzfbcSJ5MzhWGPuz/Y81rLoNhQh6eSuDojxLK64FDBUi0eSYws1y+BM
jdsrW0muW7sdWVFTyIVCtW5ULCSDuMg88cd7UrTJfU4s3YUh6110uMGuVZPva5iu
8i3+xdkG6iLLOnbIIaJUUvUuXo/0FGUvVcNFlBMf1hQ4zGU71tOULfAZ+j9J/A8+
TFsqhDVwaWuxh5FJjwUkDrRkGAH5M7vCw4d0HDn3GwoQS10/ZIJlxuWqOv3+rPrW
z1saai/8p+0u5uDyZjWBozsKB2O0/vYGEryubNJTicHqD0Vro3DUUQQd1xq4S9Dk
XZyGHw/IbMHIq7JlzzKKZ5qHHgu1gfisUxhm4+xSQQuNA3UmVlrdggQk10Ol1Y07
IcUvTEOO4L/FQhIfGs31omAIYaDUUqVDrOpHL5CjjK6XgZbkAmmLl0nI2/8xzak5
8utJT8MZ7YZxYVHfKTTRDBSM0yn22/hLe65XQ+v9klDxibtqw17FPz0E+P5Qv1Sl
RTprfUKiYcg9y3unSswrDVkJVGoflL9bjpN0zhgxzSIWy8NGKblCAjGbb58Dx4NP
I/ImOoTojEoTP6CL7yFMs3wugCAn1vPoIfnQgYMuMNIh2ucKJcAiBOnPeRsb9pdF
eeDB9PuYnn+QJH8eYiVVSjisVj0ea/cX2/UKoXMuSmx9nT/czE/iH4kqk1rPy9XB
GEy6UeThq4MWMcW5ttNxHYznSQbfDT5kFkBgWrWirw/3LQ263J1dmtVpy2Q3Zv3W
VrsBQ8V+DKv5rcQ/5dV/Pc+Fx+B/teaIkA5OfI16wfJJf3qK69z1wZfrrb8JKLJp
2nwMWiFGBPD5QGbq68kEYdjKBmTBDsbwm9Zihs5raRnihEI3JTXUqTYTPO7YUGhR
960bsQsjtElUOR8+fjkPksVzZX8BGQ9Z97HTlZ6X5sao4+EJEUyOB5vxkMm8r9ZA
KI7zFU7EVpdFu6LgIWLKo840Y2S19teLWypM3JUU4lHkskoQHrWR/l1aT1zLfYss
F/6ca6Z/50kOy5jgZstmF9PFgIlpL7EvuhDnbue8z5WFt700+G3+LlDLYLhTUzGK
XBXM9Ek31j0PmgoN2JoQYZ69VeCnZj/EV7I1ESh8tnTSCkeQ8xFshH8W1NECGFkK
jFPtsubCp6xq5+LkDawlHQLS9BjsLq31pQ+s0MJMMC85eZtKb1mGtiGP49olf0cm
GjN6Rg8ZCpO68ajbU3XK8CRwYGe84pYE1m+T1MLfx8qIjgn3I59kbb3/Pamf8jFs
vfh21KXKs5YAObXeNYtJ3yeH+hDhLzBVdtvYW7RnATHw4B5otLjMgaGUdaAjY/MB
mDHuH2mwU3Qja/De7gJdXOYM8JtmW17T3yscjyG1bh6D0enH2DQqat25gOdwrCtH
WP+I3Yq4hmKvJYuVbSTF2c3s5SnZb5/q069VPDtEABHpfSdNqz60V3ZBtQ2ludq1
FQVXmvV5wzYDC8H2koXrrPfhQTJfwMTAf4PscE/x0CQpHvbw02dBr4kZruARhuya
5iTLtS60ti7zYXt6mbpmFfQm9Zi9gTkbBZEs8gECaD+o5gqGtKQvy8+BqTFlmqxK
8i7sKn3U/pRWTrdKIcT8q+bANZBAT4g5f6n9hMLgiB1pP0KmZeYsvMWXWAaT0xzd
pSmWU+tHsdHVWKb4amujJv7KS0n6b0Ir/k1vvHaAm8J3H6cvQ1lTC8/TNYSE9y0w
Esq5o0uULHHJwvdtv7dy9QywlXmoIOQJnQ+h9Po5kl5i15gh7SOXwAu8qX5FoS5O
JGSOUePwPXb/rnfQ7bA4/xKqVhQwjgAFCoamIPsDwzZgSOkzGagosZqShoL0jX0v
Q7uTmWUOK+6jRftISzqGVkWkTEZt9tCsyM4lrPMQeIcaGyVO908REtV3D+4IgFoL
oKsbSqyfV3O0CBO4J3iil1eDmFmPpVPdL9Ss/XWcezsT+cyTvDR6394VJCdMIDSN
nZE2UmyiZUFFla4iDs6C8XOu+GBdqlHpZT6aIr6c0sCbbC8equtRHi3ok/mS22/i
GnZLqwU7UrYd6idMHlO1kGz+COlE0xR/L35rQe1hMmdvUMPtcvba/AmLkwDMsEgi
TAGmRdFPohGdqdg2LXF0cWKIfft3voHUKoiQvb1zTb8er8/c8ht5dwKJjmsmOiUt
lVdA5XD8I0HnTqXx3cVcLcaSzLSY6YhGbNuCrLxj2zQWqCkvisP3KmkFiZBZMB17
hzyBS+6cN9cQVta8WBzzxGi6sPaAWXOEJ3MKzxMWPBaHiBJqlYwhwln7TkCmnxRM
cysFNl9LBtalKw1Tcl1/A9W2rtRf/7iKXT/cUZCSGrKRNIPZRPUJML+RaztYsD8l
`pragma protect end_protected
