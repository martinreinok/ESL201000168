// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 03:52:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qjnYbEaxefbyxmw0Wl2pb2pRXDdyvSD3YPv6cTQljDElsYKiM52Akqk13I3eAF7R
zWc80d5Cf6NHrCCgZWPjh7lWC4o5XOYgmv6LaSWswf4lDvjmZDoBnQti04gXGOKd
jrn4FYr6irrsKQQen3NxoVkv27fEM55zUWXOKqANxdI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17184)
eQ+XBPO4XHQ4yow/ARZC8QIO0KRPkCAPwQkKFHXasAsS8T6tu0nEkXyi/Zp3UBG8
EvuGOZZOH37Kea0FdzTsHPZ3ieShfz6Aalwlxi0aFiiLXt5scELOVJ4xSkOVRLZN
67zJDmJBz/sTwYrxR++THPWblQHLfqyC5KQXcQozxMefzhWbfNh3R9KlED6DvZQt
oKDpb70PPt0s9pik3j3Ix16rBqiiKBrB4Wb2AlfiVn2iZSRWncJfBaSlmdrQYjnf
1m0vQ9IMf9vNe0krk4/jEO1iHTi40gGdI9bl+e1S3opMbfRbFddZURG+FezMKXQN
wJc3hbxSzzHMjR/ryzktCi99br3GfUYASEOKyMcTTsBrup59tQNlPaLNrzxjImO5
pPwektbh5wDyOlBNNEbhyeZueZYzj220I+zAkdK92ANN5vuIwJcaxe2832aNf7Il
aSlY9mCMyRU/fL2Z9ofwK5Z2naaoByJDv5hnxrx3sPEimVSm8Q4yzRQ/lxhAUGHp
7zxClCcOPIc5NyMu4rwZ3TTyEmE7kUDuV/B6pBUtqnzT6cN0oUwYI3xBGGd6jC0S
L9SB4hK16YrxXNg51e5y2Hy58QCnw3EthK5MUZqHBIRPtTMqZFvphWtDPXMesrsU
sZHeDgHDqHvy03Z1fhgNVV3pitG2nvKEOVGtLsWgJ+fCBN/AbxW7RVuTOo1tkyWu
9gr3DggTq0wBEVQLQREHMq4RUkCms2I6tRj2kBTBR8vlwr1iMjBJJWhHkYLlurMY
dCxG536Nundwm0lAPXjELnnnopXZlzoM+wChLwhuHOcbDCRkMyKnwb0jkn31dgmV
mtihAON7098p55vX/ifWjhGX24nBchZcylaLmzDLCRnQ04uHCutgPu7RtAIn8wr3
Kl+mP9How6OJ7PSdUJumbwQytLoBWU1so4NwR6sSx/R42t5WLlJRvPWBmH9VlP4r
Ekzd1tTDCTmLj8LE72s3S99bH3iUftrtzgnWiINekF5oMr3cUOiYTerEZyxsSc2x
VjhX9NnoClp3N+b68sqq/iYOy/pn5hfozL//6m82ABXfg/JfbQiyYdYf5qLJUAwa
syd04KL66H51zCFzLpXJvGGTya9q4uuuzTOMbvDSI4RoToTvuOwHLFFKof7PLb7w
0UroeNVSyDDSE758RTsZHWNB4bu5qDtNGjWJqLkBh8fcsHomZWrmw34aciVt/e62
J0EWGqap2uIQfn6TEw/PXfLLKCNDk8CNgSvziLGcyDEOaCiGAzFYSvTII/eFiifP
PGzIBsQSZjLTUKyLr/TZoHio2Sx+gNHzS0FqsFANVlpA3RR0mYbXqPtusni7hwVd
nnNm4S3qH3MUshneqmD/4rqWLxosqHIzCMdzrN1n4Mwrjor+bCfbOq83bNPbwtOC
6IThhINFL54fY1LPFFmgpf6WQ3QgJmYAdro8uyZkvUcGpEGb3YtFsM3u/wEHCofe
ZdSPqAYbMAZyV7wnrWxfQmxFH9N76ao5/0OG1rdo1FSVnpnp6lpRKDD0yFnqt3TY
rx0tlNpJGjUu2kEUir/JivLLqvTFqlHI6n+Mn8XxUwEFDI76o9rQjtmEYUYu33yG
ArQQGi7zSoGJ3qaZWhYCrIyT8++Dy2+Ubqp1+fr0G2c57Bg4+ANOa1iI6mo699Pz
rrr24KjCGAUTV9m8uAGCIwZfrcZMDInuwisZtMOnMgEU4ECHHfvUDDbp724ZkPyg
XaMVwe35SGIyK9V2O23I2IHp10nnNUjL59K8KwTIC1WyEo5Oe+iIW7V/9tv1xoiI
VRg6KO2j/HQ7dBONMtorFw9FV1mclj3K9VxMQfCcqPgxgPkQ/pxNq0+JumsZCtP7
PXcPguVs4cJuV5YLIkX+XxedRwAyo4HhSowmwR2NFpWXkiIK61N46C+CcJp5f42q
p+E+OHlmPB+t1h2BncPEluW4WNtgsFzjOKhPp9DQXYsyfRY/x6ic4lhnEWsOj9VL
g2mK9Ju0oIKSaIi6S5ayuGf6KFW2fHqlgEn+bg8+T8DVuQAWgExp+HCQqXems7+/
mpwCQ6AVtezsLL5pga2DU7e065479IdxZ0olTgOh8r85e4/J9tJx0/FMpSLVmFS9
FbADMr2ChlA01+9/Gg7PCPvhlwolapzpVDaduRgqDt57SBLdVSHfHEU6dMJiXCwQ
+NwsQRjRkN/cr2mcOXjjZ+PTx/uVCJxAkL928aLb/yfVQzo3/mhA/eQzj6lz8N9Q
hVfu3ICKxnypoWQzuqkEDayh2YuClxSUsU1FLMbetbcglqR/3Z1yevafUhyMFr6c
lWGjVBHClLrHopj/kgsz07IIBXNtkWkhXjnAvqvFQhl2n0Z27rdkrDNCobNHgEVy
mosR3wpR8kn2q58xg4N78X7kvrFGbw+Uoy7tUDD272eBlZyAQcYcwM+0QH0Q8xgW
qPZZt34iqyE+cxIr/fgIz/wWMaaLyfr+l7/e2+ItSoNHWrnAphcEh+rdwRrNC9OB
hd1OS8BuONeDw7UBR81TQXgNRwrxj90vdkoanMbR6JA3rfVVhgBSFaKZOCwTV6/7
vJy5vhxo4QWFiM+J4yp5C+zCmxM/3Hj527kmJHL9bLTTDHpF7fboN9dgYbE4LgKW
M7U1H712NKKNKeteo8/lkDPW/cIPvbGdkOaWCxLHsrZnIgjUTdUv98RFlqVcq8XZ
YwNMPAleXKX2FQepXDm0DqTPqHVhGxD5XSSHpdZKsUaZyGQTCrJnEumQlv4fyILq
5kpFmse7lQ76cASgR2r9imVXmH3pH1KKYue8/nLjeFDUSgfpLf5cbbCe57Z4edPx
U9WdJ0PW0Yxd5yDgKeTVdjPAKdsABW4l/LPPpcAXvNRw+1PS6yslPA9O3GiujLZb
LWTyNrOgsDWVbusCAWGzU5TqtW6qPwPI1rF0568ZNZpvUr4usMzOA5O1qCgBMMmh
R31+nx+WlSCyv4TIfFMFLaB8RH5xoymGhWR06NfALxBFUBYUOeCfLPdGBpQtmO0W
TzxTmRULY2ZIxLGct7ELbqm9z+PqRXkGnYCFGfdkFSUs7C4ZCKPAV+GmMxnxK9Zo
gxlBCErj5RiFdOrp3Yqt719RbgQZN6ZCXoZ/VrhfxYftz+ndqJBh4ldb9vW6GgDn
lvsjmydVKozqvup5KjogPg0oq6YCv8XeDI1UM6Qp9pLuKoDrwN/uN4l93b8Q/5gP
kSCiNg/F/f3x7+GQ69iKVwqKuUxD4hUhCJH13JYNylvQhFjdW6CQVZ17WbNvH60S
9JuGkE53bYN8SNPlbl5jF7oxI+t5OU9YvqHK01DZHOCD4TN7D7GFvvtWOfMHv1ku
dzo1EqNxtRjiRl3TL01uUJ7uxem7loUCzfQEGv5qYKuQv/+sepi3PL0flwp7dAwh
aEhTMNdS5yvfcaSebOC+vAkhOUYWs538C/XMIrdgGR0RCGtl9qtbtyl6cUE9+OyK
VsXvWVZv5L9ZLJAV/4FPispIpIiRQEy2unzd3N1p3m3Uk1ES/CKsYvST4V44zO6U
cpMzEFUAMVhnQUGdLGP24r/nmHB0vFVa1Kt496psVcUZY3EOo9c49gDYN30gRkw6
8htiXEqPgY3EB/cNWt0zxJrCCL0uBKhiX8EptXubEXHU4QxidvAPTU8aet20Tu/d
sge+8raRb4gjwDYwvt3ZCBAxVgNTXJp3QfqR9SWTgkxkDdBnqAMT9xdzEcLTW1oE
/mQdYo7BRMdxkA8cR5HPnPSUPg4bDRiKIHpZDa3Hb+UGedPoZWooxDvcFykQBw7J
Y85jVFnj2qEZStl8kwiAWyQdigtFD5Z7MIU93hg1ob9Fc6Qqmt+NTaEpBkzeoQ4n
Bsm1jWjt8FIxcZyXU289GjmZk24x9CRToBGS4l34YVJPgCzS/YBRjv/SmOoTkATh
2/ek/TSrHKIW2+Hb16SIi8jD3G94QzGNcDmbQ9b0Y8g3Db0ukD9dZU4yQcqcmPQs
VvvEAcfg0uNLunvax3hmItKsicYvCYKdJfHmmtVqcpSk/Gav1A9tAra740dgYv7f
veK/taW74TVNjIZIaKvlmgLxr8IcGasFira2ADE740aFamSu1tc7Sp0DPPUY4CD9
uxXqwfmjkEn8jka4y0dVWbikN7eccN0isLFhaccP+w9hHVbmPlSbyWvyGsKUSaEQ
Py1cYKiWgiPP/L0OZ9YvpzOblDytblguTlsGg0cFmZdVC9qDBitmm8R93G1u1xpR
s2E+3Ofa7ZQYhqQEuY+pdJAvnFJJ7n0TxN63HNP20Czg5Kjyw6Z5K8H+iTeB8i4o
Hg3F5Xip4rDCvsLxfrcbEbI33rIATu3u6PmiZmekCsjEyUd34XlX8wjSDrKEQ0y6
csQXZa619hgGzXFRdMT6952005dScTI20jlmLK+M1V2mFOHyE/LpoOaii0iTNvk9
Uut8IqsKjLbMEH7k+xn4mgapub9n4GsdGGtEt8bW6EO//C6R9M1am4OEN9aulTXO
rMRiKUkK0fzoUPDka4aWFY+Z+bL1a9fCAQVB5mddhKkfoG/F6uk0di759cPq9th5
vTnIeT8GHTBuuDKJueLDc9tKp3xEswBarCxVF/7BHcuoxFNzgMOJdX6Jb6XManoP
Mj8x14AUvzGypAVcynPNzbOiBaLLsgu0chV7YvSoLHG6EihUhOPAQaxNyukaMBlc
mbSIzQTZ+vZqDRwgdCBYM0gOZMyGwc50jqj3/0BNlbHwFrTK2c2POeKdrBpGvd8n
sm4jpSHYLQrsnpLqnk1Cu4BM7nOpi/Tm33CoiT0A73YWKx1iZuptQStpreJETriB
/GG4ce+0GdhFVLJ8J18k39i1qeUvDNnND7bjDtm7VOMnsm7ucaGojoM04hTsrfAT
Ew5Mfdjtbbpdh+hzjZ3zyPiOqDuZMrgcDhBodYvtVq0pN+/t6loLeGcD7hj9UvRZ
1kjBZSZpJNVeB0+Z/KTuGIfUrbEfRuMq/vCZ/kAw5VWi7MgSHPaE7ms//SePst76
LWTYGOVSzMA89rkCB4CaXoyleajqU8zAD8/TO9UFAGgpwhzR4NDsD5lg743boa/H
0JydReULjYmCjrnN6JVvGbokRIKNCwASiIzjgMpwEtthcTneD1qnZh7naLePjzmv
N+0en00BdrNd19IlyFQATgRo+oLICY58COPTq6sNdXGVD7PROdnIySdIimdhF5KE
vCp4u8t66F9ddZkqruap+RK8aBjLzaYlK00+3LCk1VBv9c3oGcth4Q7zcdH44y0a
Cv52DwwaB/z96PTUBS4PkiAp8JEVzXDGyNDQOePGdce5dpX5MND886lw6SGGkMQv
VJp5vaTU0Tccuf+WJNZ90uFeF5z6rmmllBGaPEZXq6MqBGf8CDyzOT9rEByZpLb5
hG/1YMEXsodm5bUhp/udFtx9bh18GyAMYypu54iWVkgkEN9qwnbwEciMztyMEurO
KjRxkuQam+f04r8QiKuWQQtU858jHH+zSTf3Kght3EpnUu6LNuZADd2c8WeuztU/
gwH85yeh2DcHvwkR8AxH9XXVPnHoupui82439SFPbRT0kwxL5utQcZPrn1K4j0Ae
Q9eoCaaBfISitSfLyqLVuLLUmP3AnHv2Im5luiH9FAxGuFBNlPk/pfwKiCLbSHkY
ZfcppkBXsKL+kWMrgM78Z6Vgrq+dGw7cgQxZxkMplmx/mM0KsDGPAiwXRt1k1zGa
mDbfag5ZMMVTc+5XQ659lw2Di9mwWC2CwRPzIFFIrtcnXs1L8JJtL8NKD5DAZ3kb
p09p9SBGxBFLY/0/KfIpiBgsSd30PmDWUNJLJOKw2iGhp0Y0lcVi6MHBzbi+9ydJ
MGuyQM2jTK+IeEaLZDVrNdHZ33kDfrW5d/khFPBLcxYaP76y9jd8gEpze9LGfcOa
3M5nTTd689FVITIhEGlZShNJU2yRYBnWzAHXOWT0Ig9u9Qo6WdIt49yIrIJNlp27
zv9eAk+fpMe3+TzUcvfd5Qq8NS6ycjnYafuD7G2CD+JUyzIxI7Qq0cxXXfoFWoQv
OSlPAvXcyv+8iGRYLHpHaewT1zrHcv6Y+/cFhATYKYLwNwA5U0+ZvptoEaBTHE1/
MAWshyxo8yDFo6KNm7jjrVVXfkmmMuNgZQY9SdV7jdLMhMg95rbjUOXH5YQfda6t
ftO166kinQtRsHEnkcm4xHp6upoVdoa9Kffecgq/or2D5W0bzq8tIMQd34jMcXCJ
OhCPdkdQ0llboVmlYmLzjiJL5rwriZc3Nqko3V+PLq9x6vxoiHC3Fkr6PXtjNp49
GvInHFEajpFSn19CkaHB2YbRCLEaWSXxAK+2jJNp5K8yqUii91MNAebe8DmBLf1o
fHsi5d71mEoDwJLv0u9jVRGZMiwM8KQXF5WdtFhcb8jYWvZLAMQaTJKyr6R4l4wL
bNe7F3ZC/yoyUWH3qitAuB++wBK2zCdK5DS/Sd8ja14gICa6MwOlB+Lu7oXAxBBg
xckAjkfdRWDZkdLgVm6GHBOXi8lx4J7hGGedL/pspZFPuD3Bq/ycOLkuZUonItsp
Z05kyT9D4rh9IqbcgvWaRNQw3VA3mAeZSw3oPfXe3DBlqq8p+1KZpwU6yqfePxZ3
bbwyMpFBwSCS/zqWbXNrDRUhMFtxZqdYskeOQngv9mHlHi1jJ7+BdSNGVLmoiU+a
cIurrZTtLnb4LOPp6F7Dj5fx+PEgwkw9jWtb9eNZzQvQwJjMksCopXufFfEei2WQ
T6LCCvvbojA1rWb2b4PYiVmIZ2bUekFu24uzMU5AE/MqD5EAt8ZukM79HUY05MQp
RT47V26ulgnFQvgwsufdb12mDD7+cFiaQjo1Ndkd0H3PMkRcLfiPmGbRTqALP8Gw
/7i489V96Nc6rNzNim6eNIkrNrhRBLSbVeNOzPbAyIXvV6aLEHryUFM6uKxpqMTc
Cnf/B0qNQWDXvg33xeo26H5RYwSAJSLrldJxJlUkmeefI0jSsAAXQ+SENRc4iUhM
jXFQQzfUkzFW4v69lq2d+cf4478MWOuhp8NLuMuXiDBNmsizbsx3ZQTEqU+dXxab
KZ55eoaQq4tskRQ+SpxlA6n1ipgzc9zsGJbCq2t0RgMwWTTt3oXrlmjd7MxjK5QW
8yFzJMEn8P8ki4EFXzk+3VncvozEdP8dPrV0q4abQvI8sI6e/aWP+x1H3T5s3c4h
gCQQjC6q2R9p4N7It0NRTRMyw/p4Fow+rojMS4s3MEHEfGQ+ONFszShos5mBXTaA
qTcGOkx5N4xizu8OMbJ9St1AgCkPapP2fh/yeb4HEa30Ic935FLu6//G2rlwGrFF
kWivTwKlIjxPnDDaaClzJb+Hfy3aZzaw9bpTosS2+aSBMw4CbCv1WUONgxmM63RX
pkaURmd4gkwBEkkENDLqi1gZeLyJWP5JN8MXloCwRBCTVqwYFh6iKgm9/RvmRrvf
4pVGzsrgLSSD07TinEwIC+zzgsPEj7XolhGrOIYD6OwCipLCiU8l4jcFqlAkxOXM
bqto+M2XWe0P31FXrtJxdjjCZZZYomnM/MI7kCABXzp/OWkpi8TtkosFmmVvmm+u
0MotoDErTk358BqVuLM6uWGGpFAEhgllg7nw9hag9zEbJ3QAr5fQALRlNm030Lls
WNCEbKsrsN7LLEFDBwue3k7yZjegVV57oFLmIpucnfMmfwuNqhcgKxxuJrw3l1ka
FAH827YO4AoKfYfuywQnlO+itPTgVa9DUcY+WIjAg/95TxvMBMMJH3MHy1zQUxKJ
u7yEKMzslZWkh9nAWLZ6Kklrcs2LhfEX69woLuAdPGdL/uppucH01ad7g9jprkJL
4aXwBcLSTPEUkzIo16j2SniwIvcm05rGBeX0wyZwK4IMyeD3cXSpX/BbXkh7DBmT
Faa+rR6sqC4gAVBxoBIQi4F5hvwru2WwZ8YeWU2ugbxn7t2mOU8k3SPJL2Xl9EWg
HPuw+J9fVYqBBMvXCFxBMOgBiVKk9MxfEr3dAoKEhsPe123kMMaMEZAVKMHaCKSG
qlAEmuHG9lw9Zv0peAIFaCxKbIuL7HUmKT0n0LgR8aHrbfFLL6UI0a4TpfHH9CEM
ecS9y6Cej1096qlYH9hdAZZv9Ulav9QTRhyNYYg8jL8STqxWZ8/sN6aF92WVi0ma
IrIBwPoQWJSNvHrURoKYTq+z2TRDwO4oFZ/xCAneHwHaVEbFjkGKU/4e4IRaDYHE
G/cQN7eVOVYuug44ZtjqdOrFbv+XFGKwwNaZ/NrxYXbDned+GVBK3+OYxE8SYkRn
LEi0rpCPI+4lnKYbUeYZqYbUD86EVmZOaZ2Mn0Rsm2mlndx0eLYLVZssO3hz9Mnw
JAjkt+LlcbFD2biXEiBgcqYou+hTK3x6RUKynv3aTj8BC+UdtnR6H7yYyZucwExO
JcB/gkQh/sBoDeMBMaoQS0G+xQv1T/7hCxC+L1otfMivMnNIS2QQMcxBoghbDcjy
PgfEf/XGdkGOhISbR8bqC/zBH9UarhkjBjjhePQFfaSWoHiCtpV7pb2lRzXTSjOR
8Q0U/Nayg0+BL4MAZn0wyjGDYFdfGm5bSWOe51mEIDvl+xelbQiWbpOp+D6dVHXi
SgN6vDa5AubG2GgN6hNX8e76StKebLH5q9sNTF1WkBgEYNLad98j3h1+fdUCe54u
fa7qJtJFe56b2i30cn0kiabpOBWFNmUkpjg59VnE2V+fiTK2V7CB+dMuTK2RZL7B
vY1aOPEn2K/hXTVKp9vn4zdri9p/2yJiYj9KDZxU/nI0VXTnWdsSMWJxhBiY5P53
TQZOEt9sM/49vMNbUmL8YW7q/Jm3NiAPJxQggYLmoVDMsexCc3gxYAOZim4UMFqr
ShWrWcFQaPUQKE3wVAKz5WfSo2Ot49Qsng6ULydRSmFetdL/NyY1km7TK2hIpVS8
B3pk1VZIDH4sauRA+dCnD3hjIgiK5x9lKHt7vsx3lnSRPKaBEw+7VZIYCdydONsw
rXgnfKPjkJlY7dtoGUdWjqGbMipwulVKqoQYmLrUwPVzHjXE2iWZzVE9pJKUbzn+
e46AUceStdAkMJY28muWM97BZgoyQXv1ERgKa+Y3P0KV5R5VQtOGLck2rQiQuHgQ
96s6KvcfCZaPgCcfXqVcsdOywIdklzB7KMslCOmpfQRJmXJAtMtdx3LD5TiCrk1k
sBF6x8l2IBFLQvH9gbSRBOBIaME7tUkf56QJDIo7if3azhdbpJeaf5D7esxD4yCG
MeR7/XjsM2IYZLIzEgs1C4jeGJk1IpTldp5T3phsa407+EQPpM5iOUaShgbb1FT1
ejnQmgF/olfnib8MdqnlAPcaq8pxovOHZ9+E7P8atDtXDDGWhDXYRTHoN2CX86GE
9D+JlXBfzbvyqSEMi76r9gKLQcUAg54yjZRM4ia6IoDoYWHYSCloTG163YbSsx5J
uQJJ1BOzHHufsieOBY7unqEZCD9ZUPOn/t3MdtBnSNt2R/CD6Nsah0dh9l4yXMqr
az8t8lUPeVuTcYpgNvS1r5gdH6rD4dQcRukyR3hLxhfDlVl9wV9xbLqqR9Y1ZA4P
LcICuJypyKZoUtqTvGqg3Avyz8+k4Y/0yBQRH31ch9xhcGRWCdk+Ku9Osn0inprc
rCC/bAepkvaTvIR/mHb89zRXysflVo/6iDgUeApKHJzmY2t6pZJQTncMoz5hDNiZ
3LQGfesJopAtROpgCMw6fbeeDN5htYXrgbQjqx8bZ7CsUVEquLnWZOaqQtmW2I9s
xqfIRQrasVd9oF5fLrSw4YGPhcBpP9YjsYhtCfGG2tyuMA/Sfmf4sH8cMCMMnL4r
OEr3Cdzemg4we81QP7vK+NgFwvE66TH5CRpH/oO2RdtefX5EpXruJcmRofmjU1lD
7h50pspWZ+3417XOycY+FuIEz5JWzyNtyPx+JPmNyx557ibpiDobAzr4UskB+M+E
wQZB73tir1jVCBLS4Hw7u7sie1XKO7UevZ2QKEcvMjZHRSJ/5eEPlVNTdX0yVXtD
2ZQe9ii5gxeJJECZ6dJwnu65vlhxda+Bl1NN3LXpVtKC1weJW+evK4ibUeguzWG6
GfZGQ0FNPcpbMrrShqr1/+6YLMjsN7gnEQMU9Co6aWs6zQtjmvNAtDQzasKvBwkl
q2l/12EN24VRo0W1CyxFzb9HbL6veB4qquk0CgGBBYw6pX4iJ/LqQOGArCjI4kp6
/qY0zM++KOvA7AgOImD0K2sYnUZ0jnWh6t9cA8SaWhfDOu7ijAMP2+rSzMpiCo0D
AI5NAxA418k0+fpmhwH78/nLuQ8MnZ0FZ6GKVhaBP6YTnOdbZhsITK5YWnL5Smyj
kwOktxr0G7viv1hby0djLNfFa3ZJ6jMot1laDFIdcqtWFG/YVuX22hhIQLz0+UqR
oAzXbLmBexFYu328zObw3OR42NnRApPeQl5H5vVVigw1T0yvSF6SV3dxtBS0vtHv
jVdaIlYCAODapWCLxit9ACI+AsS9rp1SH+2jAt98Kmv5vFzsKXsPd1i8Wszeq+Pl
khQVfJ5nHrf8AuXnp9o7i/lUdOgGNUnSTF3eov9FO77bK69dDOwLSL20dchsbB1R
iRm8MI01McYCepQ3/2saToC7boeunURV8abcbRsNb1Tn3/eLn6CZ7Jc9RE9r64U1
95ZGz+CLuPrXXWrKOTWMX5Aia0MnZ2Ah4OOhSlDY5LQ/ZtLhJPSiqQXc87V3Bv4l
lRb7M06RXRjyediCmZI++wQcJ88fYNKvve26AaJIoEBechQCjNcnBDwyKqV7AQo2
XCp3g6t7O14OEB6kL/vL2+YNPV1hYf2bh+y5ufivjCwMgqbNxyRbnuGXfvOvjo2j
0W3fsAtEFAtQhkIo3GfQMWgp2VrXuMwwLrbM0UQ5GGzzWh81CzllYrFYT0PriJab
JIFhX84ZZEzAOmTZnAGNCUyjEtvaSfDYivuoHnu0fl6kBo3oYUR4xt9/bn/LaEQV
ooCHbIK0XB0nDFy5bybxxlzUS5M/TN1kivLSTC1sQLFgUXgvIMdAS5sKvKoroQzk
aT3cF/6f7sZgCktm0/1EMnXmZcuv13unvtIWjhjeo64ymuuBuhDwiznnpkLLi9/H
TTbtsOH+mX2FZ5jl4jnec46dDzfaE28UelGC8U1Nir+a7R1P6kbkfi38iissc8eF
WYxYEi07TqjkBRDkG/1tDczDR0ZKbAPbAeBExD04YR4bRvjOiMV/tO/ZgiWbqbg4
1FO4eiW0bfjyVJPx8eGqavDL2wTRkeEUNMq36RIzspGRM7//qYNCsp1tymaE7hep
rMH5Avxu93CHmZ/SyUAspMRpDdJFcqxr708ijsmRofMO7195iBg9GBjPA/31j3kr
e3x0SKMFZA4IUsKVMcLn7aN9+v/1Tfculn+1Z4kuSF/v/d9+k4K3dtIxIxgXIAVs
Ip/HJKAb6ABzv7S3CPv6uWQq1pV2ytwtWrjrpNMlilO6Er2oiKdSULIF5wWOHlh9
jSH5xwpElEfJKNVGseGbAiLSDaTYGIZUm1xnZnncuczibXZmKAuJ7SnPoW9XZl5V
uX9cIuXE8IHhsxTe3LYgMEPOf8doaK4KJbM0v71GX19TyIfVHSGrF9aCD5BEAoss
Iz/PddcyJ2I92BtU9DjsIXRfJpablLJV7sIczrAs5rFxdeDfbbrySB+H64EqolH3
/q6/noNvyZaFZtMPHCSMOrwlidXNr1eexFB9OEp4sdH2YR34RCTmKU1R+8ckUWy5
4EQiCG7A//6cA/ceOhulq2cS+jDy9ovqxFSX8RyyICSRs/HjvQJFc/Z7OAM4R8if
AH4npctCM7HB6e18GCJCj5HYbxsRS1XqeMSVMADV6XubkaRB+VfWyXQCnuDnDGXj
cBrcsL+lwaeHdPi5VTIl+355h+q4rWV/a3lwGrOr6kuI8yqyfhlbt2t9W2nI1SjL
G21XrY9j0M4ELG7RCh9w+3zodJjGtOFQixpRiuXuNLQ947flzAjtWzh7waSPRV6A
tcyi4giZMsNKOLC7ZIGYEBeb0OsfC1s72ilWK36hClTAkA6qO//7kdB/Qjj1P2hY
30AWk00kDwXMnYdMveMXs536UC2NzlCMifmBZVrPKZorU7I5KJRiq0p0iLPUW3Ht
XWwmq7HaSDsaFev7eUcAqKmtBuP1mjCuDRks9qi2+IEyRbOxHdg10lE3eEzS1t0g
ka2YkiohBWm9bk+fMhR2hraZ/3dN6H+LtOdGGLtcebYU4whgMPqvRZrLs+lMkOzX
siYfywQaXaXeY3gnmBvJcdc3cCWDG3XT0XK1bAhl/dcGrjyv9jTymMSZsJl9Ht7E
ibXAT4/jQ1jjiQq5QjJJnAJAyjGrY7l3mkhpYQbk4980ioW1DqK1QvoLiUKBLysr
DMWIVCtrHvIlKZciHSGu5NHHFqV0QOK5Cuj9FgoHHNopyVfxnjS6zwJA154p2a8Q
ZkZVG12/9Oabb0I1hvvMTG6bJmhyHq59IJJv41oWh1SiW6HyFv4T377NkQrA4SpV
I3uUXvsEaR2mMRF1sim1OZe0rrUHDFG+5CqtAb8u4xUBaxtEcrnfSCwG7xV8mydD
Ei951cb9jOGXRbRe1KSs/eZR8KrOg6LZN1mOf+kVn97MgDh96HGFg1bt4BOzfsYg
iPmE4+r/oZhnXVitPYSG+R81mSBbMYYuR83fdsg5n6wgJpFJ9fy++UsEo1/CUeYN
27Az1nwFS6Abc3wzf8geYz7Tyv5FRPXVkRGEHWm59brt24KucdmyGFLF5ZkMlnYN
j2XgDIG/s0BeK0jrKX8jvkMb19wEEcF19t3If7SLV9v8JA6VkEwE0DEWYJWV+ptm
uZnYaJ/7f51W8VXSNcbLHFbuymE/y4MRwTvFrXsnyApAouBEnnVnuN8Iqtu62sCf
pwomE7yuR2dZQ8knOR7fZEuhNqd2uJ+CWxIFg4+/N9xDr3rt4c0uAzrmAQc2fRVK
ZJFLPerNoHD90LSsF5/TtfP9qQZxLqvtsW2+I6YvuDv21XhGrMFmWgpumdrEJeCu
PXrWQt5yn3FmKaLlYi4HvsJXaCB7rdsQmTSXpklG+ukC5iIbcjAQu5uGef/Cvffl
tmjaJSlVsfGk+KTOih1Hnsv1IiWDoBC9YkMyh3O16doZP3tUd4gk3KUdf+Z91tD/
oz+ihx/Pl3GOZXVmGCJeBQKgaINhxvkOlUp4vFHaE2QgLzMxULcCdohjiu7Jbjd9
O6LDacyXsSpKtpoBpXCT1YQYnPPUBlwDaWr7xgaYvP9Hm9xp/mczFHN2cxfAat2H
Bpe+0DhKw/8VNc8h/b4Gvdi74YquWh7cbHW99pc6xy4hzQ/YV/01YFE8AX0xq0B2
XqvjqaDwXiqnQJeoyHTdLZj8Y8Nj8AcgV+cs5SBGpabAJBuls1l79hC8MSOnL25U
muFlyZM10XYLg/eLtFBNsbh7CNZmL1opKk6LlAFfOWqamMXMbjsoDTiUj4bA68h5
rT86YpnFH5dKwDYyBYn3rOxhbsdPgP9RWCRpyYzRZLjmiBRD2/2OR8mpsed3JDuX
P4jDESVbjuSFGXA87Q0sFYB7Tv2zbBAKmyf5dSb5tSB6J99/e5x9zcZ3iUdWukDl
MJRtydIEKOR0AcdGTuOi3Dpu5ea/qqGBQvdMYCTEXx/Fs6trusnae3GaMeyx5tkW
yBNNBw8XJ3rc7bVQ6ZTUfIWQcFQUfzqEeUIF4T2BQlafU8aqX6pwvzbhZg9GfYRl
VEdS3hYR+wzBVVmW3m+uaMLaaWS+2jXrDjNl+19xPNyaIU5ZVSNR47FFkP7zEFjS
AUBF2s91wtIB/ZIFUs59qAeqzMdOvsRhJ3tO35BaxiRngTTGFtn+q8e229YKvVJ0
fez6Lp56c6+yYr14elWFrf4VVSOn30oiFV0BhQOkjyZhChvLaAAQZ5y6QMyYMi5H
alJOhyohyWTHe8izqSI2P6DfJ8a2VOI/0Nh1ph807LQi7M+HBIgk8CMRiJ7LHUAJ
e8TK3qFMM+FqMzpQQnMFp6C46s5j4OOjmFjk9zsKOrNfJ8n7T7ndLZLn10wlK/e+
ql8a9MUSJXm5RG5RufvpAKcMvBy/AEdvW+oHjjLnYEZcxspsyfJhlspFfcBIHSjO
fC8drRK2jxfxLfM4BPbNHhWuiCm2PCtrfY2KroZ4+kubTE94SSu2nA+gmNztltvT
rSZ6O/UXgv5IxwPME2t5ghMp0ygKEkIRzqjYKr0v7BIWwEVsD3xoTe8Ediy34Fqx
JOSfG6oG0oNyfU1ixQj3unvdHl01Oh7lY2Hoov6d3YONRxB4CDAPPFKU2tRjO6vc
W23Cg/u8if02nfuk6eYS/JFcxGM0loEiy+t1UBwLvmTLFYe39VhbBcoWegMefokk
+JX5yyJgNBX+T0WJaXyOqrGiWOGceRHxbhcjyKKkVoy/zhKSfeM4sF8augL19Ccp
hbWnWqC4zKuPfUsu7cx1IijBBgUBXXW+Do+03zQaJOH7rDsfMhZySsIeT9Zz8N1B
apPSWleNLhLvprqX6WsL4otfApAA1AWVnL1hf71bGIZlbrc0xMTJOQUc0Kz54+8p
lzgpUwYEEuSioaujDbqc8gNjceqhdrMb+3S0rG2n+o+JEl3Fp7nz44Y5gDGcrgR5
7zi4wnDJdiYc95J0IQuU2F6erWxkK+notK9LjJ8jK5Pe+0Lf0bH43BCMDxGbNOnO
neKlbfgE9kzCgbPmBYB7IFF6N3Ara0MZOqXwF8oN2/8OjcOYDshVUKQgWZslECkC
4kBsqzMzVDWy0D1O/6cxJklY00QFE1PwDiFvuy6hTEa25ycjdDPfxQdaCURHxBTi
HShzIJSrUDZ/QrZ5tA9jtZ0e0EG9Pdu8KksmcEzdNdKW1Thz3Yia8rRXw2yGOslh
fmnqmKt1kZRfEY9/tEfTDzm0+EJDiWBg6rTKCTBdeoQxra1+uOFXp8cuX83LrT1B
vcd9ryHTp7Uow6hp7mmPp+iX+IIHiBdiEt2kCcxX27WNO01fHN4nTtgI8cgcqEpR
V/ouwpNj0zRxBFNci6h50PfHh3W7+KALGwq0X4WEn/zaEmkkvZ8ojGj70URUjsDh
zWkI7xN/Nw7Sc6wiwOgdgP18J7DrRAjcg1rRCNO7W8YAMvbxqVhf61mUWGQA98O+
ti02n6xdMi7Va5qmRgBMfZXNsmch00Y32uWcHhAYeOFgd8tPnj5/SLX1ZFlC1Wrq
k3SxMAUPXBrMSsaiiIFFLTvCDspLEUyFplSThRwUd52T1x/vePwZbgVoY1xAf3tf
2JluhP58UciFH1IqIpLNZsdQfqM50wjB8T9zaaXIpNHLVYGZxC4egxREpBnWjraw
Ltteavqp5XnKS3wjYvrhHM3RVx9PDuSc17EYlgmxLAn6gy2bE6KVnsab+hm3Bo5I
mOdbtlT7ocHOE08TzWsMvaoRl0R1Sa2Yqt4JApuGR6z52ff2hfTdvBXBzLAycHdl
tzyBm6iFLo2rAhAc8q7JspNJT7VAZ+LYB9xJfxHdMDiMIEdA9njZsDy13/D4nFTc
brxkVIRwDnJDfySR1dF4klWYWHJ2IbPu1yeeRfFixcTdyyXKRiqgrIwCjGkRPfFV
z86yldhTn+t3rdbNCZJwfsuz93xQLa1szUuzU7TQhVWzr0nUyNo1MCt9e0gnivhr
UfEk54hWYB+iyXd6uOBxEaAZTlsVQiykElxp2GFK/yL0pWWDcQIGMYSBgBPdBI9x
N/tmcRCqbJrUCDDm4o6+iM1pBxhmOE8+j+CEhtbgBIr0njVp2C+cEex2v/Y6gMNQ
0ILhDfbUa2GdnXO8FRVo71gC61tLYPm/e0lBQ0vXteUnIcvijrVUn5g/rDW8367P
YQ1qAmiTohll/gs4OogjPUBtq4ymHXI5FZLZwMrxlXqunxjzaWpj9fQxGTlWClcb
Y91NVYnhRqnC1SR5s20Ld0FoiFCneZWsnZ/zKhIfSyR4kX1RXEw8uKua1fIVTIsz
M30TwelKNJO+s5qRBvWU92VvYzVcQ9PjmHpPOlwW8RMbiLL/Lco3MDVju7W041jh
uklSGtN2gZTRtBi1RCmRmB0phBDpA+hwSfumwdegysLIozTcKIutjjOEjctmpJGf
f+1X99UQuDhWuvoko7ZwrMMucl2tElDtczt/xfe7GwNt6vtLryB/D5CtSzwNnUYX
SFR/jKbUuZuMd6ahJCpfvToCcWNOhmtIRknn/jQg2XcbnIr92jYwuaKM9jijskVj
gzpONmhl/m7k0XxVFb4LZxxjgnh506RmyfM7Addal8R2++yRABCKBRKB6gczRsEe
A6IYgsXuiWa6v0QnrkX3dgCJXEYcj2ffBI4jRQF0nATgsEGYeR/j3vQNYfgEttJX
XxAje5IcZBK+hSzstCIsSEiYEEl+MyqWVIfCtAPRNU5d/f0sTrTUKwz9BCy3P0wD
9Ifq2u6FtB4R2Qyz8BToV2fykVm4w56PtmUmSIWA4OJBduxjZJ80mXVA4gjfpYMK
B9sag9/Un82U3BmtttD/j314Jnd0MWvstWZnnxwXVGoqH5Dgg7g2SDEDeDxw2+RQ
w0vXCEG+CTHJNICHDyrONwsLQu/Qqdj81sEb19YnzAEKnt97vom2yBcButvBTIa7
x8OL71aKeEiZfurMetwdsz3Ehg9Q6EMUnpoU1eJDAP98fnqfSvd7LCxN49PkwpRe
t6ACp6Q+dvJqDkZ+Vk5bj/SR9W2xrf56jKhjpAIAfYLZo7WaofTJIp42smRE/3Ho
qo0gtp7xz7wvMIpGc+GgwFyqp0N6y9IAnargqxLBPOo8Lt+wITOpKkQSll2JMQ3y
XYlXsEKYadnNKQgZrU8wNsKjopzCZOawVmhVLuOEIQh2qoCCppLS2liXdGu/TW2Y
p4HZU7/BrNSTXvLgDFm2E8gm8hQsXKCN3VwYcY2JlntEEfBBeYBCuoo6Qx7ziI4g
et1ARvNaLSo+7q7DjAlK2czF3Z4sbkYpV30zxcp95FGToSQ3xqX2Tv91Z2t25fRY
EZclauElC0dRmKS2lTV8K++ScIYg3A0MzelskUs14TyFkAKuwO8VYR5/vCdSv6sJ
sErLn/O/h22U+qnDRK/MBeCZZxpUasLQil15Oi7BSA8i4KFkpv1VHbdkz6C3TrHR
+hyJIpc25YvanRZpHmZk7oXwC9uNe5wScCROzF5GjbsXK+qNfS4lf40UoNTeJMGE
vv6i58/whAEpiIRPrksyDucKdk9jSWOq3gQOLHAhIBQKsk/ohcrHGydm/WEI/IlD
hb7lUN081Cl9AkZJkQPzChCl+vojR3DzwPpIefuxBUr+uHb9sXKCaraeK5hSE+ev
gnScJV6we4BedFoFPPAZCQhVnvhwMIpLucNZxROfigr/Wx2SmcNqFrTkaZ8mtxRB
p+3fX66U6RAz0T1CFv+aBwETINrmcceson8bpY7a3XqLqTfDl87lGB+iKFggTNef
Hxuosl1vxpw201vszwNpJboYMQJvcJvPUXgHV4YKYql4CXQDjScjlu0duUj5b7Ty
HWcGwiRndYCiYMBY9aTnW7EofB4KTYxvs1eOeXBEUSxK1QCfmMdCnTREM2UYV4eR
/6q6bDp9CevK0ZMZRGsSwSPrkfPtWuiUeWamTFZ2D8kRx/kE4BAOwO7ssw5N+NJy
jotNGiEq4AwrnmpWs9R4D8CvN/yMCaSTP1t7n6JQSsDKyrgdhSyFpD70AKkfZ1Jc
f4/5aKPoVBDwbkCzRrbiRJi9Vu4JWSwZXXXEsMDsj07dyGxXXn5+eB0h61EE3bqN
rQD/nt4LXgHLwvBJJymSo1tLanotmASpbFUzLE8CEIZ0q4EezCsD8lsR0NAvmOL4
ZPwmhidSt/HmVcQF+GV2Kpsw2/Fo4CRax6B8g/nudfcHfNS8topW1vWKkvUyOtsu
tORe17rv01rCiMqknXarMGwjrBTTvGWhnGDFPudXp+G/wB/rzzIXuFj521Vpi5hq
slsP1sPMFWs/mKuCUdP00IR8i2MAIMV/UM048bzN/B3yWU2tTfEgfcD5nUE8sjb4
gruxZZvuqsVUMVRsmHgjldb6T6fwpeKsMPPls62r+mP9b8tFMvyPwmKGsiYUgVcd
A2yEHNHNzNhuBD3fvA2pweMIi9t66vmeF+UfkLRbK89KiOy0RqDu5q+F3QL+uQwc
NrRFziOshuxcYR8dZ+f1JQHtnFrHjqHqN282ZZ1nFRaMofJwHfl73D6W0ar9RVLJ
mtDhjeKdxuwlBofu9mSVn6bz3JfwdrAh7Til36ChdIq5L0Hiqbu0a3zjyeqFGcaQ
0BO/2EcmDnJBgxvzwGwLdjoAOdqdU31iORog+RGo6MwBA0XzaPE3C18Qk51VhpuQ
Ex+PjYl7pJouCfTubG1jdwAvYMa1uOhdD5bl+hVMcytROgA8/G+DprgWM55EFWXC
7nh2O48JrzJFaMyLK1kiPmmrTzzDfeg2q1R48xBwTRCX3grhkmMrmrh7qF6gyFQf
zrqyBwguPyLqKp/F0xC1UjHx/k31kyiKKR1WadeNtv7KCCLdr67s2SJ04KdJB+xV
gSPremLDbgAwamJ9rYUDD32E9Y8PlObkAQ/LxrBLaA+G7tlPlTEfSQteYz0wkoFu
q5ERf0zOBnaDKyuxasDgcaaTrDW2RWd////8GDwRit/Qu6VE8/e0N+5muhytLiW9
XgMkBHw15iIanhksDf9KH3wrR+zkk3J7D1fh+vdNVliAKssimjoh2gGkRN7c/STX
35oTL9L4q0GOqZqKPj84VWh1gztZjvZehiLEymF3qOKW7LZyISMjsrCBiA7FOLY3
VPURROODiK9eic4KM8hbxW3IitKUcHGTt2ZiPxsLa4QVm6JgnrgG0F4k/QkWctGv
96rrHLXtNNJ18E1A4UVogirWquA4h8AhEfoa6gYSL543m5z4PnFErcy5/ycoGObc
ZVTroBnuqQpZUURG10to9VjdEXRDvRGuTJ6UMo4zPBgJ/bEr7c67tPmhUmyy5qli
OvgB2kY+g88y4pzGnQ/U33t3sXvlJszerhaBkN3vCdUFYLbIXiiw4S293NTldvcC
RupG6vWNFvVcnR2mlvJBD4T1NZG8dUPMas5hqclJkppdCSFas69sWnvdb77BgJZ0
iJIJOQ8gRVy5an8SKmU0SZGNoLCUC1dnWVGgI2185f7dzkMxR2AneXc5e538eDL2
ZU+QRMRd6huCd0xkeGDeeRKqgdTEhdLhHgX6YuHEHUw03eqmBQtrjoJtHSN/toKL
Yunj4iLtYU1ELSLhmG60/wajza3ZULkOZIfdfJdSC6GPEhGONcFUpAyUEcD3hhug
tRm24lZLZnMaz8iEoqXhtFIUTHzF9t7piUdMyH0ov2wByxcgAOeGW628+vU76ftx
bCnTmdRsC7nVqzzH4fEXh274wo14kYdVHeEowoKu3siIq5DnEXWVMYCGwoHKUalB
+SU48xnauotqlH8CjJ3P+dazGCtswvCNnm4BHkJ5C5ezRUa56yzg6l55qgcJpUR6
YJC34mhwTlphtT7QhJumj1QOEMysqF64v2RxXtf1ZgyRcz8Z3cmC0mSj06XiNu53
VkqhbRuzCu3AhFi6mTi7YGSmGnrXKjxuJMYZftTO6TFcOlrdtVfWtHL7G23vFifQ
88OzudDxY7YFu7LdJYgS8WkHFIprtKvswx37fFNSgz1H7yzQpc43e6J8sAEaTuEa
XDjyNdhzSwKHlxtFjyZ7Wi67SCYW996t1pzVw1Um0/ezVu/Bix3n7PZirytPBhNL
5M2aL/Y4EWSaFeTbnt8COiRH3G3cu9DRE4FMTxYfIXfPJvqknSJLbulWfGjsqS6V
gtMSSvSjL0HCWUWLoz8a18irFAm4UsxS+PEKJMRWdNZFFGiNVpg8VxqS71RgCvcD
wIuU1BI49YACzKzrGAqJ202o8Fe+eANshTixKqYh2LKMvawH9Kp1NnEQ0m9pGnAk
VWw9RKOxlaFC2zjymuLfTYfTLrmGxhjpTf4RUka+/gER8qc2uTLPDeDfxMDWV/r2
PutCG5JHsh6+PEv4DqlAIwcp7/OSNLE/kYj5zUF4csKMQ4GxgWgG8cwNDTGHQJky
NQ63DOIL7bAOyjCrId7oAJufskEU5hxwoO79PaOG8zolOZKGFTs9oMsfPdiFx/bZ
hAzVXm4rIGqOX2WYKvwF30PLXzcAIlFAWVSIGAlwNdYvdMXlQ23TY2HQokMgiUBg
S3TeS0JpI0VJD5+KfmfDNYs3QAlT2xY13goLMbj4yLjVUemOKB/Pk7/7cv5gkDQk
9zkVUkT+4uZobKzCMCsu6Uno63tPBBgJeBwyw9NlOC1wS0m5bfPMua/rXLxio+jz
TktFX94joHJ2TC/lIFXIuXCucRKs0VdKis+2XArTr/TyGi5sdUfgtJ+6HXff2+pz
p46AvjqNqQPZWxaGcMs7hCcNC38Z3lTuJIt10rgiJg8r6HOKtySDf/ZzgSDQ97AO
OsML+UhhUsaeLUiqFf16/T3RlMwjyJhbaLYcz3R8NqjKAgBSw7ZQjtBLYIui03nE
ksq+CXu7oqcd/RU2f2vTrzx9ULb0rrMWsjeuM2TjKpBuLXmMEzs80jvJw3g3Ce0D
KDmCDve23miZ4vKu9/6aV9Vtc0dk2UOTC6v2o1RgGe74SSfFIbb2jo+z3p+wspT7
f6rWBkbaN8ClEooBdAgnT8EE9A3fHpqzLWgnJItPOyzGF+FJ5AaVQ6VsmkMQfF/G
fmt5zEPAGfw+TOl0VaWPB0Sq/HbsKIRISsJQ062YoTJImfiNmMulQag7HKsaCtkI
qc5uIKbGCm23nxVa3eafWZXjOcGgGQsNG6P/373ZE3Li2Rf0X6FXvcpRbajo3Yt/
sZhBFkIWvl45AYP3xutXLJrBAKF8zsg8UrYjoWnUI2Ryh29JTUjKWfy7GnG6mY/G
GjkNCKBQcJ5ErxbcTFiCH+La/Yzka/ZjaDJcoXF65CMTqGFWlD+G+EazGelU84k8
tC1ee646EdJddIvH4X4/a7H8BhS4QC9D9HciXN8c7JTERA0dXW+Q+R611ZziWRfM
J6CZY4hoGZPD27Iy97hRO85zzNOIFFynerv+AZymirm70DMo6UQJ0f12U5zgHpqj
b9Br9DOowUdgvQ26cbeSc/mimCNEgqW/qxFbScREKjObNTl/sLmlp85xTI0lpcC1
Up12MuQsBBxy2fecAs+CgZyxvU+Tbwkj4/tRLKH8/+rZOoehP1/WoMtyz2c5rIlH
OZy+EJWmj+W/6fVm1Tyyh9qNWRCkq4aRM37ywtC7uEnJ1YQIvDpTCGjs5t9lSAfD
0hPv61XCn1uOp+DYCxsIlLxRmXgaFJ9M6+VgA6NgeY6RpYw+r051xQNaauODC9FL
zz8X6DklMWtu15F5QFZipI/EATdVSBIEpgqsf3rSfvjEspAVuiZdkjh9YsqMyBDm
T2VYEQASgaL+47KYPpRN1QzQZQCB5Jn7H1W/XNFk2vkZ+lYrnBhDgf7wAIpqnIYd
V4Uh4wyqNlmXPzN4Y/uCpau+fby7xrnUeeqf77a/1BuqRvBKydM/ieqBgZj07i72
GFNCWyavUmhD0hexLRjsNq06uZomeWkSyGlumsLM/mNhRvhpCoUaXAIrcx7n4YDR
nirFIQ3AuvL7pUKHbcxxM9pQyfTVx6Lg7OpyMu8ueeujSzro6FrIzsac1mr+VtbC
oxhFgWfseXr1OGixnQwJcbjh7NURDnKiq0gwyi4aUeegWC+1SBbJOjUXtBwAeUqi
PUEdfZTmTENjvY0ZfPq2H+HbdD9Z/t5sjNqsfeLpAV7tdkIXxFkjwO2uIpSgMgX4
rWIFU6gR0oOUV8OUIuyA7tOvQgNb8a2jiqvvpfzmD9TlRSHp2SQBL+1QoG6wU4rW
E8loGnoiqEnCPUyolaCAtSj/rdyp0xyUk+n52zr1zyZOGNuvTIRttRM3LOHL/7dR
QZ912//C7OHIb7r/EDeEfrIOcv8atjC1MqcnmUKQll6ZJOTIamGc8O18PF8JNjtJ
3CnSAKiZVExYyLVZeOhLd9w4Tm9JtPHBZMF6OE6+vE81GbBKQeCHPTmfuKSg2Dho
ibunVq9eioAP7tkoO3SVu1Tv9WXgOAZhZPIqyoIaRg8HIIiIvggp1d8YYNh2mh0a
a+g84J+YKKpNffajrZOMUr+yn895MnVUXM1TkZ8s4rFuSQu2o1914F24xHeA5qtq
tlb7gPhPaJ8kaM6+qrCovdb2D4w5s7u4MAx8HA0mZ76tzML2IW6X0qE8uLfVbefn
Ls+fvKiYeMzhbDDnM77E9t1U/XSeY3tg/mTkrPADtiVThovCPB6Qnw4j/XLRD5qx
OgRfQEnP4bJwwvARRzSF5eQiHTjW/WELU+pyXAhwMIRtd2jZV1Fr/E2AI1DJTtAr
mkl2UlMZbABqu4DxQyIM4em/a+wy9aQJN2Mhcfi1cPcBsxZV03y4uvY1pFtFT+la
QZ6T8tgMtNwT+frPUZ0HE8YMpLWzIg+tc+mYMNRjU4y5nkTYJTllEGHH6nJNt5Hv
t6cFBUbI9YsNd/5S9i9LX9sTiOUB3I7dLyEOuwxpUXNoYDhd4DJ0RDIUjbPn0p1P
OBANvhSHQFmijpaJlzKxTQWRf1RQLmfgDM0QKDMpKs4pLCV7gmnOpNphGEc45bdA
9RF2nTesyaRe86SxOwlEXBMnhyskhS9cMxWy2TJ/w6OXJWnO6ir3g5M06Yq/HpnS
8k5oByAyGInf8zPcqAXb45+ziGhylUfy2UO98lxqhb6NmrSngslQMh8CjasvhF0D
5zPfCNBEn7tvoyI7qx0KQT1uIDyQOOkO2Lr5Yd51LGmxX0Hc/bmEG+E5YzmWMkJv
WOCtJ0giVSHAShv4f0ZmDCzslUyFW0OHBLDFcLXWf5NqkYpTy3drOIPWK8eXaiq6
KFG8/QtKabw49iMT+hVOw8CRcSWhi7Fi4LuTtPlsXUgaiQkQSeKsjXCcLaj8lfh7
`pragma protect end_protected
