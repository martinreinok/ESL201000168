// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
UIIPA5hgViMXUUu3CkcpNGozUtftc6HOv0swJ20Qcky1uWzAnxWGk5z7ieE77oYV
lqCdvr3s6DuI0gn1t1Fs5VU6ozSlrA+XYba43fjZViaCX+9oQZeYO5PUKlqf+nRf
dVjxQAE1xPxrrd4dCcwG07iWhqkk07vvUyHGzGltTgJzBRlCFbln/Q==
//pragma protect end_key_block
//pragma protect digest_block
p5JRbMYSFykkADgrStbeaHTdvHE=
//pragma protect end_digest_block
//pragma protect data_block
Ai/BAkouDWevyLW1Q+RTvBisyNtbYQbQiKhs4FjyDuNe419awtB4+Os/LjGOAOUA
6OOurzjt9g1h7ez4fmBm5I1SD4UmFhOxJejfKRX2GfWuMOaHSP8vi3VVJjWJ4IFS
CvioGlU5eUOQY05ejp1LvdExgcZECFAwReBYCmV3hAJvlZYuh+DDyfbieWGDE7h+
nE3Tf5k3z5sX58zAYZRAAqm8BVRb4QtfFBQMlOiwVI8nx1zEPV3KyWqHuqkUeD+5
5w9SVi/tw4nU7e9KcBQeEYrfXuig0BLie++m/7zrVent8zGgvad1QkijIiAGN8Ah
g65ET9p0F8A+cTORzd7LCXIwxR7+reMG7guPOWKnVRfNA8elTJIed7pzcKZPZqF4
dd1OppCh+sK4vi3/6gsAXzPdtw7FFEQ4B97HN8rZozUOKqGK/zY6oJ5dsGnHrf0n
vNbExCODaD8JzBvXtBt3Zw7OFl0RB4fcag59YPrHSIgrfVvt4qHGQirNDwuMHdwG
2LArqhzarTVVctxGPdwbfgFt2OHksqrLZvewm4jr+Xh3TLztBz/qVo4mbDQEIAVS
4IS0lqt5BX0o+BxZGG9/eWCTqdpaGj7MTXKY4rX+oxv7WWBOuODxxZ6YSlwIcY1E
byHS64X5yhuC4M9PUopVdQ6UxUMOE29PJOt+HHDSgn6o6GGnp2qAnQfkS8Pgft4F
K/xnO0rMsbvmp0gd0b5V3MwP6/uk6Wd+1lNyyv/Y/JOlI5jZnB8X9daH6R1RRkYA
r+oRfoWnrMeEvXem/gk10YgAKggAAdm7qDt8oky0JHojH4qISHLiPcxbR7jylW4N
So+OPHNJNhmMfb71xOE4qcShIng/l1+xFI2e6xDVd14Vx/sQXUOG05NgBXf2t43v
NoF2hBDZXn9mskcc+k59AYPqAr8tDGBfkiscJWZA1w/as3YzKB12MOhM/W9CU7tL
WwISUr1wXYww0A1Zh+wE/7AFdFMQ3cTw6dluXMLbqd2KO7/QldHy3uJ7G/KtAiu3
v9VRrt2cCfLg8OfSpRsksljjH/zKVbx6+HFfqBz43k1nURb7uR9Z4lrQ5lMeTiL2
tx3QGO5LeiH56fIOSrjzTdbiD+aJT8UnAgI2maUW5osdcYyeCS4x6MF4VucpTDK2
moicV4ncvzciqx6K6SfcJJ+Xtc2iUQvEQxxKMrszYAnQ1OVw6rUADH8PcpYBjdvE
H/oXnowGYnppR87KCM0qBSaLdUO9MUyLq1Cyjaz2zcX4JwJguusVwQ07BomRV21Z
JbjtzAb0v1Z6BmTBkgNWBqWtySFFpO2tqM1+LcagKbgzKx5qT4cIosdGVpW50J+V
wFR5Q7haPTIsH7kvM+Z7MLw+FTpowijxof2+wOQFkw2x6TMgRJe4QS7MKnwEEwHH
cgWkzF9UxGnEkxa+f50h6vm95BHIxUYWgTRPS1h3w98OuNUng3UcpskWxxvHOfHY
nocVmgt/ZvjYHa8IwxDFY/oTCdzUQPbzHLCprktYi7FfbFhqPAXeVrXRZK/tKS8Q
yEOpk43yQSk0nYwB8frAOT298V17q5K+ul+RuPuTyTuAqBnzVwdq0VF6oUz+Y6t8
6bT9KMyt2RHi7B1M0iXNy1dnfwoKhJ+UuAqV6Urgb5r37+aOU4ngkMIOx75uQzkv
VHruYgeWDqPob2hfht9G2ujWSnIYY9vIcn2rzKMC4RxJF5W1+PSKJX8kC0tv+0jC
Kj5v+yiLN+5bK+Ze5diP8kO53NRIJG4DTHC+U2Av44to5bCFuo4O/k/0rA8UT6hB
GemMCfWI5y1vydkd6fVubHPU7uHAeDfNjssPMgHo7263jbuLhY0XVAnEnAG3v7u3
jj7szd5UwVswwZdEEes5kh8tbjdKDQVQlgMDgKAsFq4RcriocaczGDZKRTop/oSY
+OJICENyWf995Bio2If/gyrGLJ0t4gmxIh/g75EzijAMk3yS1NTQJxqvIBnYse0l
b6BIUlVRb0WTRVRuTfDyLIe+rR8uqND7rFRL6fe+B7s8bJHdlFqoCQ2ct6f01Gkn
wv3+aqqzKT1+VIxH7isShu++X6TH94P0rG8/a9HtNjZp2G2GzNJu4IJzeNJ7wZdi
VxOEHJajAcnDqdUUbgEf+Qe3Rk++DdhhHwGCRN9TiS9E+yR8WZoulyWpQvxU9ssg
cB1jpNYNMyQLXkqNOGnSfb4cbFD+K+h2YjBV1zuML3Xx0z1Rj3IGRqSPE5+fIWAH
7m4w1RJ0O5AfM5k5QJWCLNwm7659px1IW44A9IZ7dR4dBedgN/GFvABVfhQD2jg+
i7WwXdvMzaaE9541Aalhex++assxply+tmlcdBBq1O5pBIxYW7MzRFu0SMEKtWcL
Lq94YXe8bBq3W17hy5iRDSwKLRrgl/i9DnM9RSQd4Dc/3s297r8/q1K8I6RPYKVA
x+sBP+TRRz9u2QDrEddP7Ng8tNg0g2DgTR9cowto9jtrtHj1t+G3VuOXu1BDVvN2
AHXshOw6eK8OtkRwPxuqT1JvjtChnhE+syuvDwOSKUNgAW3oiK+LsDZfqvJUqNTC
6/csGE/TkuvZ54IxO7fAzhIbw90kNjN9oB7rwYnY2gdrhqP81T4DtNf5wO5tkr3E
+kcSql/tHlpm1kVfLF5+MohV7aiPDUuLsFP13DG3Vtux904IbUXtudgud7QOY26I
kI6/IyVIrcYRtVEEpaDIonWeJVJ97ME6DftrpaWu4WEi0pp61AdxBXIzuAQ3SqIe
yn4UibRaqbjWUlvtAeRNrhA8wA54KIq0e+EV3dP+WM9G4OBxFDUeMjamXvSkc8iG
VMMSojBnZKyMLPra9uc8zN0pHyoHEpmTzVz0MdBrEIRPeJebwNyL8ICHKWiUw4RF
TbVbNsVdDIsunuJZTyJUusMPKyaX+hwFq45jrSkHbiYWVUhmabzQvzgefoWHPfJO
FQSH0enJ5xXMCSXioCMq/nf/ebzHT3qjB7207PZ6+kuXWmg03jH8a/UvrQItoFyi
QCxe1IBt1kLRMPE1noZPdWW6vcARtr5IpJnkY7mdoHjQXXLwLvVRPmQbIWTdrwar
7u9t5dJYFghobD+5SZUihUFvvnDh6gf0teZfXwW9Y4oXMXDx3WG4e5/TJ4womzTt
nNb9DRe3hURzx6eIXn3PjLXL+NGS76RCXfDEXdAaNIxFcT1m6SMu7TvjpCSo7Icq
WQ6gNGjDXuwNSIG1a9waOqpzx6MtrBlIt6hr46Bc6LnTIH00FhliVizLAOgmP6QC
DmCQMXTzP2Oz51Ajti9TEK3l8x4G+n8NOvFIA3UktGdAx3vfYdvuaevtGuILuEmA
dPYyLeOMCTyPOYULJHh44dX8VFX0QUogBiGz96hKEjrMdvXdRbxwJaIuIa8qsgeJ
psn7S3Umdv56ELIO1uxllOtX2A3/Mw9A+njTINLIBHdfyDzsdUO8It7eg4BwaO6N
Ub/qw0O5u7ZxsiisBFI0HBb1SNlWz4Kp9XgPqUxtCL9c2G5J7sGHLK6H3vX+RY61
W6zn2AZqogdFh1A3N/l1PtUDw1RV5f1k+l1G+SBLBrQZbfhU88Rngozko06SKCU9
8URrF4PvBzBccBUq4Lq8TkcEiwiSaDmpCQ+j6E8jS5rOv+1QQiu6H/uQ9unqxUpQ
FECFIK3EPp9QgVt7tWO933S7EdTRONUGIkPMD6QBrL8YglZtVqBt9DAWykXyya6I
bzElVvx+mRbXJvt0sQEbj4TFkJWcA/3CNGQh41LGy11Am7Cq318UEK+bAuId5ptO
rcH3r0guiSW4uN2vvmU4E6VFjtHirV3iVN/5v911wVbYTmAE9/yJq0Z1+F/rYxCk
IVWngo3ioNzqrsiGkj/B9iQB3SLXv1N6ZV/nmoqQ+vb+Z8OZLNscOmjcY8YcRWIR
TVx8fNimSF3ENxPdOg4KlLwEkVim/RScbBdpStf5qRdC9/ImBtk1HruEgzoCdu+x
nsDTiUn2hG9UqMxTRDsb1fBqIcI8PSNB8scYHDp2U8XZK4gTBxOT4h57VLi4eO7H
UEdFx2oDkdtsPhw4a/yk5LP/dh1IZB65Qmb2zfWaS/FavZzW0UH0YJZpRcJAH9g1
ZKSfUTygnLzVNwclin6HgW0Aj1mEJqfTA4/6hLSrVGRA8725r6tfeONzTEeyKKEK
sAGb8zAt8JjAzYjM1kbB1SmXjLg3T0s5GEfcdVno+BRIxPFJzdykJD+Taq+2YFcR
Af/ca/ovd8bSLs3vHPVkJ1IOhK1DZd5C0xM+/UvPuZhk40jJQmvQXihprxnOedee
2GKZXohw4wFRNFoBAmf8VZvEJVssw6il4xgMU3YTsqmEqPlX/J1R+/13X3pA08BA
wCvMZhsvr6fAlDD6M38isIgtlBlc5bybo8sWgZ9ryQF7YubRE8VmqqmLtPOLeilk
XZGOiRQ8Rxp/c+HxRgmh7aO37aUQjpGT5fZ8U9j0Q9YVjKE6iDYKf/3DjPiJHhBQ
GAJ29GSIm9FdTOAoyGL5P+BPHX9CBe4Tcbsm0LUetERtIySa7/S+J+t3srinmXUZ
98wOonHYZc2i3UvWEO3WPFdaocRB9aZi0dYWrzrN0UOnISMC3SU14cdN61rlM7FM
oF64MJm9t9Kd4YftUhwrgXjxT4LSmu10qZut46jmbca4gySfnw8Xr8WcKWle3zSf
Y35q0+DbPGlYFq13iQ+Ag4VVPhEkopfmJBoUT6ntixzQ9VN9Bk3yBrogl7EbZZHa
mMDVmkN9/HjvvH35w7r6hPCN0d8liS0imrxaSkLpF9wT2KhzEqxk7ny2iZFrz/Ku
nh0zMJ4rGRHvild+BQXeiZhPuRxhWXiiWIqy9eySIOFynRE2JS3p4N7OsU+hEwn3
wsiIHzzJU9+OjsU7sNBW9LBiIQxO4jAw9A13SG52RKRzvhlMSgV4nZ9fgMADJLS0
OvDbh5PvWLXr5I0/Rdw8dR7UahMMQ9L7jEmNPW78TYudTwJJH9CUJobRPMTA+Hbg
WfdjavDijnA05xtnd5COYh4qxbaH07jpfMtDeQWOAjbylzKkfbW+1o9pwsBFWc1U
2DME9WsWZYQrpHG2icix0HgApg76GmM9D4/H5gmt1wXzWJcVCpey4rClgMHvxG6U
W3pY4lAGsq/qqJbnMRdw6xLUG91GcUmPxLFOGVCZtv7zk05hwBbPmlC+iPJ4B/6/
ASPWMrknvwhiSaLsd4Hxo7+Ao5LIaNgL+bchEL82WC7cxYtqerwdEN1p+h4GHM8R
DqitsWrymZeD+qCYQJfYPjSuJkw5MRD61Gfxrb72o8ywcRr4vTJ40JAZ2/MM2Pll
O0SKbjk44mGiNvgw0twBmsfRPR/Q7fMF1dhmdV3np4um+bKZoXFzEi5FvWipmUd6
4wkug4NaGIPiGN2Dq6tWiOQKw3QyusqvSzHd1Qfafqs0o1DUJ6j3MyA2iJ+RoTxQ
BfGdFBzkpfjddMHIx8rsakXFtqEhPkMDwkmm8tQv4d0cENdVsZhGiwi300hue6jN
9o6VmsQjtBtGhNMHW9aZC0MV9uQ+bVer766fWTBUwQbZiAu7eC7j/5PGNlzmQJMu
A4IYn+SSYkvWS25H3gIVr/MSgEWzM57glX09LmgLfBZ2QtsMu/Zk/Q8mSTH7EWQe
/xmBJd4luWxocMP4KWDUs8DdiP/AORFQWOo9rZHZ/11CofTqBDS9wLOOJ90QW3da
q/gbkAb5v0uRczCjY2YZIZCZtv8GfIoNn0BX7G9tvDx5EnDEqLrxuTkQ+z13nXHe
Bh/DBeRTKlSDo/jSKlMpN/3WeanV59lfRABQvyBZXG6QVubKwLHMtvFbFHhUm0qH
pvZvoZr1Rz317PQaYbl8W/uFB9hyVlN3NBik1xvgqb1av3Vhw8zD442QJKP5ryhW
dWkwJzCFgtGPC/vgDQjNTZ7D2h30rvqjLJMv/lWMbCSilLjE6qOOfcnRtZdyDRaP
pHaSM+3SRxfo18JGV8e6kPxd9Co//+9Lizwi2d3aFHWAMyq/oQjXIJ5CnBY5FT1Y
xRbci6nSbGO/BhB0I2Je8iKkuj5TOK1z5BFvpjSw+hGtZ6eVuWLsT91S2FkdmA9d
uK7CtpQbidAFaWW9HcHVn2Jh7+6rziK0nwDdNgEiXkbrheUsIbZnXKJ8iuCZNg6o
QWs9aTmYK9lSWpP6rb0AhCBA/T+WMCDcL39N0RfxUR/O9uVhA110Wx0IOUxw8Nys
XfskHOrjIPS8swzIqqPVfF2PqD0800K1szCJXPx8A1E4pr+hb+dDSdS34TgAKHm/
YzyETVkY0FlzKwE++5s9OsaeDrtkIaAuX1AJ/PMN7thP33LZjff/ibLoJ765qNfx
3qIaxRTH6wIdOZHPOu6TlqfMH69ktib8V1KDzri8gsES5CZhC1POt5UWKZvdiFtb
qY+6EA25kGKjGZLeHRKzA9OP83KQadN42h8IJSAgb/UwqcXvwwy29I579MkTvjMG
CuZtq6mD1Fpn/u/eYHJTj0TevWUhGlVNFQsaplj14/etiIBatqcqhc7JtIyo4B9K
MlgFMOz0G1W9zOuTUmk0hawJjFHfbMwy9On6LjkoFSUq/MKKwwfcjxgB80Vj4UFT
879CDSXvDrGVJ5GA7DbPyMtYLRerX0kNrMF5AB5PBRhO+MTJHfCujFnLCYAaPrg7
+/4GQaOiJSsS0fo78zLSRtda881CfouFYHgBxQXU71bZTJVIAtlPxDMnlARo5c3N
zkQwm83KNhPml6wJsyTWJta7f+l72BCc5yf7FFsooCbPz5fDm+3h5T4AfYAoY405
mKmWhGhHF2L4OK4q1kdKn82NrofTmOVCRZh8KGzIev8wLX3g4WJwHnCbwL9dCTYY
8IETGYIQYdhZT7XQWqfxc26FoOWbWlj3qdBykYxGqewBo85teLDoe8Kb7XFz8WL/
raKecBp3ljKjcFB0tf187rqz/G7pZq8vWPKIKtTTV4MfEAaxII/nVPZvlaVQtitV
GNVdh37u6gNiQnXIkIRDxerc45AC6BLdYEdmizJ+TJoakhw1/h6LDIkxnp1eFOKC
LDa/I/hPjzlRJnVKR9Ir0rfrmL6M8hxdxCPw7nABmVXXcaXG8UmkKKEFGGy+UFfR
qOQWUqVN4kg9Gb+y+y7TijjdG/mxoV3vT2cPFqhnbzA5+iBYHBZzAFD2pHf8TGAE
lcHaAH+3JjUzee9LHsSkCutvl7hg9LBOIuomPK5/7RdrYqvGbeOROreYvffmx2RH
Pcvh9ELrKauhD9BObJgstnXydd/qc0QKA5iKLhkY7lfFWDBuNGJO9RYj/DOVqZxK
7XLwyRVCGZL8DiEguQA+DfLNAgKPgGN5v6acgwkodLcvcRUtEjF5r/ta5YSCC4JL
qf9CCHrY9oejAVjWBLExG/VP1qVpaWpUWvu5p4r7v4s3V50FOOuwGOi2/SzQFTf+
5nDzvXkInA/PyR1QetYCoaEETydDNSnlm1eqqmw7asa8Y8Itvj0/5hHvsDmsQKBg
psR4Iwd9K3cYiCQyybtWeznJKAJZ5BxR36Pea7lfNkljnkf4QDtICKMm5INBmgOZ
JwKuJbqqoQGrZK7j6j/BL4s61mRym+wfoDTiKjh7isZYbhPp5E+B0nEsiRSx7YUf
qi89/55eKSQNLeGU7/iu3Pl19DR/Ui1aFzl8oZnoYN0yYbIH3JCjCM/Mt+DOqWzL
CbtMf0XM3DdJLfVTzFjgEVNsF4E2v5mLT8z460B4ZsZuOaLb08uCHgfy7OPTH/yL
T8wa0CTSa7Y9LGoBsO1RuE4HvBkgd4Q47xNikchbJLYfj9v+A+vwSf/pXSqqgPhr
75pz/fXoTt3ZPU0TrWCfxQ4FcoyX3QFEVDISy0q7tiHnF49QoghCzUPCJUttr+tF
cveqlrsZPxPA58nm+lp/R6FSMqONO3MaZUnAPpAlQB8Z4KCuGulm84uswD/+7tHb
ZApAza0npuil9TTMjhR3CCh4P9kcINEqUJNrKOSetSkcJfdSHqzBbrdJ5mCOLToX
Rnu+oGIZ2QhvaoH660qs7zh+69DwONyv2xNvDGWAu8CZoKQhgMHK+Ah5/fg8jbN/
5DgMgw2R/89uzyvzrIW1d8kLkz08XUti9lpKb9sQobcETq9K7OP0SbdSAWI7q2CB
A9wDkngHii7x9EnfIzf2sAXioLtL4ztpYV0c/g+9/DAScef4wx8Y404kgYc+1ol3
jiS/DN/hHU58xvjKQdktTfIkkzOj0zTSTW0I10pZjMOdK389MQ9s2wT7GTKDZQSe
vlV0A0loZxqYcxV4AlFaLn4HRz03kXCfJgM9FKZLctnaR4j+rh2NSD/E4FgMniQd
AoD4oG9Y87sX2QMi6ckXRzLouJ+Z4UbTGlhnc2xMQ5tCmPFrFmeiDL+1VXO1/XOb
L3Y+6y80TM4S9+vN3Ot0jivt4jtMp/jA2CA2mZ1yAsbZZ8GdQ148ObiXiLTzDm5J
HPAjfXVPGSEt88opWsRPTP8rUQJha4IGEL6FD0TEYSKnqIziH6HBNwiiQTdUtKUB
nAVcXbac0hhhB5FpWDQ2pV0Zt+aR0Gd+HbodOStKXncZXT9epCLg8UOuEjpZzCzo
uZFFhgEbHQB1llqbvsM4DJSXFOMiAn1jJmennFIh/8BMgcrV3nSVuA+tq6k8fuUp
wKWaayVQKISTdDDA3E3fAkeeNX8+8m5BoA85y8kUPaWczqaDTDnwPbbpXe3Rx+rJ
Wb3fn9la+frTOoofXDKq/DOu6D9GO8WDwAIox/LNEnXbGT7AQTjTvAa3pvaMTPM9
z9KTOrNHkKRWbEcRF4p9pw1Zo2ZLkSpS5pYev/kuQLvOdawArZOQ8lBFxKhbk1G9
2KULgrWseS7LLFZGKcKiU99Lrr+RedS+IYlLboy4eQv3bgoOwaZstD61OhcNvIKD
Tw0PMrhpjZ/aOOoynnOV/SGCEyB3x6MGnQERIUDcodPRBL1QUFBleLSoIObddlvD
qBT4WqpZGncmXV/2oIggPFUBjQ37qNJnYh15/nTmqgJrNgMfVRWOq9kuXyG87Ax+
8vg8wmqPQ3glCASumb2h+eR3jK4k6/rgn0eFIPUL31w+/uWegVxkr/uMOXZby/xo
Ou69a3J/rhbWIyQCcgyNt24RDwM5wPWX1qCxugpievC4JhLNCssyNLKtC0lAqUtu
GeZb7YUDYlaKpgau3X9+S6j4mnHdx8kv0BCIj862v6+xUg8AAcw657j02qMwU/gS
kZnRRdOfEwX2hlJCAWQTciUG9LzH4tGy1hBY79+fxcJrjNQGohB6ze9hog0XQfJ9
beKDRoHLSJLJYtTr28D9C6Pkh8S3C4mMhs6XcAKM6jrb1f+D8eF80/cbQ7gJDmGp
WlSsufFUELz9WfOr4F5wCO/8N1kbjP1FzZgeDp8CN3wTrcvkupgy35579ra3IUk7
iqEdn5jOsDW1pHqjgtpx06qFwexVJKYWocKetTO8nUOEC+Z7BLgTpvK/52MT3+qW
PD6RHIJPO2koRtByQwBagp9AK/pvdizPFHSg8CUsZ7K11D6v/+dYvHcBrWUg62HE
1b5T5h15bxAMTK7NyhzWcxCBL8cGUeZ5k2GqVOBEjJfnalOej7XnZ07BzX35k5dV
rbfTYipFhhidky9a3rrWgykqPKclbTSAICRvdfyAlCe/0qEHsi+/jPsnX/9CBnf8
iS3Qx8/A0+mI7+8TEn9ySAmSThX4Z3jS+SbOu3Q9hwwikt4NE33tkDi02VxqhEd+
9cSyBvWfSYFIctSOIRmaHxfhkhKgSc2JxMgNIjWfEdUsLz/YhJzznDRJq2j5Yckq
X57gfqdGfyB8TLzbt2Q/edDkHq5RKSNMK0QRJSUHD7sWSjVOV/SPZRmRJMUSPo+z
IMxMdwMtML5EL0yOAgo8mMIGmwhL9dn+5B7txH1+2zOt7eu0pco7tcrLuEgLbR2s
4w8QhW0ZBKVxT9IbBPPnqJyymxJp6z0AuIqYlMxWJKfjql0u77puLFVJ/mvjFSwZ
ladyBaaygv220H62UyUBMHOQGdktysCAFsOwppcI0LxjP+GhWrjpYPIR3EhI7Tlt
gRChQl+h51eNzkwDK7keeVA51Gp/ccXMGTR1NpPjNP5yb0nGaJilUpzJ766MTf3T
w/iRFZQ2RtpcvrXBTz7XEqlVQe7plK/aOon7QV47oVHm3c98WuwWs0hWvvU7mCKo
X+q1B9nZ2eTys+MTMo+ocHU2x3LGPgjuR9dBNy9RMlHEc0d7Ut7We60LH4Eig914
z5saNe3DB0/pPHsMlyduMLiWVapgJX3YTBninXOU8gBZVQhcQ18A8PNaOVbbqU5K
iJ7pgQS0Edg9J0VqeFK6ofM4kWKI6ReTsPzEj9REug9dQkeDOuM7/TCIkDBo5/Gx
I73hFgNcJ8dX4aYZ0SMSuuKIVHWjDfGb+lVpVelcHu1k1xsghb5S3JVyLHCUzuzz
MECDI1U+cDG0SumkJuf0YeYqP1EFbRQB1s2rWYMEYwbR6GBFrjqZyLMMBYhP+y8/
GhEWz7b+nuon614tDJ7UrInco/AxXFHscnW13IsAjzeF973zcPzL61wqWUELCjPC
DN7UB1qmHfy8feJlydgdCU5hitmH1dmT07HqXUGRbpDpgPKo4Oz5tnz7i9nDS2Kc
E6yUKW4NiuzNqAr3j/Ag02fHAoHAwVqoZarzD5472IJ7MBGEwL8YZCjLIWcVuM1U
+OsUQdN1twhUw0rVvcYYXqvRii+dfN51PL6Jc6I1SMFlDgnvobPJKdgxTxtvPNjp
xOiOtnEYeb22oCriKEZwqHYjF5izhGdWACJc75tX894WyPLyJFdTKb+ot/JbSv9g
o+djNqgaIjZL16SuZI1Nn7MVFdoK065mWdf5+N8JeHRUlFNX0T6jkeEL4g6leNIe
pGj9QxFtpl8vTtpRRUhtfNCp1EYDNqbyMyodHkckT1fIMR8N/7Ah8SBBrIyLjHCG
k83PsFPlnFjKqsi7aOiu57ye0Z7REJR6rOErOwb3Hci4xV2jCWE7a43+RMCljeDH
t4SVV7WmJ1z1u9r6idMOexOdIRhFFdUt69O3Nbn86+R3kLM8OVqY7KXt18WSVhqE
7j0AD0Scwk3ZuZQhWpOJh/oPG7UEbbXPpreKGRDCWmK6ppj/zoRnSyNGdMVUUbBD
dyZRVwrpmWLdEuQEv9DCSpG+DcNDxD0T0+I+t51joy3/+VRzr7kyUoVPrV/8sUg8
tXI+i1NGXKcjILaYXvxHbob547QHZC4w241BoguGi1bRcdqbR2tVdSW3CFffg5/+
DAkV30+E/1h1lfbdSExI9C+X3dpSxEgjNBz1/aDp/mkYNVCJ2CHw/6R/Txt5q/3T
Aui6mP2l+VKogdPc0GNGARr5F1K9kZx2iRFBO9IBLalKcR0QbCByUMnfhHNjdvmA
6njY58ZbbnmcJIYqYjpZ8ouwRJaz0BCcjX5t5qwu31U1adiXxywyzKalglDnL1Hq
3YbsoD/z65rhf6F7/xJl4eSBJ6rAMVKNE4CEPMASLlD5Xf7q6MTZJ4+Wa3unaFys
3AruWiBxU8pfwcM24taNRd2xeDK9ymKj+oL6rRKdl8aFGNfl8ycHzQhGzlqq+xdH
SNgwXzqAEtj6+mngcH9KrGMqugEV8rhRQmVoEUoqoyUjz7s3ET+dDnfWkYz8aRGy
sjFanf6EGhDqQdepVwsbO0KxKbD3MyeIMkqaCb6hmXmMWzDYG/128nsLD/jOhE/M
QY4pd4CC06BVrAV9XP6lCQLp/sVrSSUQuAuUXqeZsKeAlouU4jfvmUVTfjZGJi/f
HbL1RtlJtgwi6s0jLPa0fqyNTgK+DEBcgMlHziEdgVj8rUOlRl3LMngKhqb2gOyb
b2QjRotXFScVhpH0I+5hEYPM+AmEwSHcXaFsW7EcobZNDdnaxajmVfJZzqTFt3y7
TJo9YEgGN2iIw+rVrCN+uojanYYJal2xd+A0zuv/qI4T+J2xFhRiv1rsg7sYFwJn
Y8WAGgMzAh8d7bO3XWV4F5JR3iPoKkQ9pmz2QMeKfjek7PfDHnFHqfAKA+jBhLa8
NPpzo7npJeK/aOIUjy0oR+f44ZELpThJFIEomwk+IrpIflnOQ4C68spI1PWYPa/W
VZ8723/sbMGEOntzn67A3u3aF0PCcTHvWEAJF2AOxLwDqL7UpP5OF7sysP98x65I
bKdd+4H/o7JtZyKrKlk6oLH2mjuE5rL2pXEYzvItYqxtS9V71j/LkcBHT5QP2+AJ
zk3Xsek/TJiJ3dtJZR2N1jcMuiZDlPIFLJt3hEDixFvKUmj2HalBs21NgCgmcfJl
elpFUAufN4FHTSjJDULOb+ePG/AlItyguOof53bJYMXTBauO2FdgXavTIsNei3Fe
nEPYJomRkzAa1XtMJ9Na/eOGh6HDhe5F62MDKq5fDvlRLvRp1HDdPVpSdmSTxsbU
onxEEsieuMGkKJw9U652yqGHEhSy/u5zarnZfRQWo+Vq005h7ve3JgDKoHI0qYM/
Yyz2gDzuHN603OR6/J5WjYa30addzAel/rEnqsMmh6ckvQboFD8VacPzddLZmnvV
Qcqz8H9RRYR4Q4wMN2nytjqx3S1zxn8SEacWda5CN1IJxXCmuQUVYAsnTaNFSxUY
TJrpcMc47dR+cER6K3guO/CGjpfUvo1P3mxf54EZsUW/o2Qd7U9SY/UXVwxQqOev
lJM0M7CU0C0Lt5Z0OTLRAMb5TexnzI8I02aUlNFsu8KhSPPlpiaKz6ZUiU5Yjpw+
c8M4paF8yFO6xqkgl6HglRDzOHDK+nQoTKniGYHdGhBnLlVhO4N6L0SmDBmnvTT1
1OSsLdPrS/CFGGLmgdYVMZWZI8OTeRZVjUukegkzzi9hHzgxU/vcXeB1/4/DqhuV
0zfQBo4R91Ce2CY5eseirgfzHOE2Ljl3YV3JRlMOZLCpu+RnV3VXYOfzQ1Xr0T+U
RKmcdx6oUsSv5lrc8W1n8/YCNIgCK0gS6sg1xUptDuDQT2iAxlsArPHKPRTWydKX
ikungxMNa1mrp4euylPdPL4o3pOa4VG278LCR8JPtlGODzAsSpWajeCyviXr5exK
b6rjudBzj9PQz327NhD7Zm+92J8imSdK52qcSbsjH4atNwnAU846sHeJRnI88c/f
qQ4pVRotYaP5CduJhxHAQc9DLQhyjbkFQnyu+RyhW41EkdTPzwSv0Bl5cb/j7JfI
CV0J7MMMJc0p2vioLMOvoDQda3EmOr6Vq+OaccJMiMTI00OKWhdPfU8HBl23SHQ5
01vEdqCpUvGnUGOqgaf26/7ZFt6ACySeFFNUcxCCmFqf7g49RyVOwSUQGL5D5BE7
2jw/cNFbFtFmgAheEQcJGIYr3/zTG9sVQ/gCfmb0Lc/I4l3Pw8NHjtCH5kcdxBpo
GrRbptTxaPDIObiBpZrr8tuieSoaqRopaUJPI6jrQs+CTz+uCoDHgZRE0SLgaiJB
bYneX6qyBD9M3b1kRfGyBMjgjN91TTvf/rtysuKjCKKKFXp3TqMXFroBW3EgJ9//
D7KLOvxWhERIk61shMuEKuPQhE0XFWQPVZ2B2BECFIXLzyX+4MIVMEU94dJQooV9
WmyfpCVJlxi4SPmCr3zI+uquzYbMnaaG7N1Y/m38kCNxVJLzazgZX+60V2rMCXeK
wxkN2b9+ycU6PHruONzbvPbEVFQuDLtFe6FTU67lslULRKKhvSwpyIh4XQKmtE+M
lzeY/fiOm+9gsEB33TYg78qWy9Qux2/Y0SdAyP9FBNKh+uBV36ZQ1caXokt0VZHv
dH+aMox3Ukh8DpeMHbci7itjKJz+DjHOhzGYbi74J/KbwA2UaKQGSUK3r9TaRsKn
oVLJYOcvcEuDpQgjeIOzgwvBgl7L3mp468rADl57AHryLtRL0RFSfjRsYqndDybj
/dsQPR8Ak48pCfQV0adS4+kgpYWPqwl01Isp/0AMoSVVMddkmvc7R/1Lrf3XlwW/
zHl9JU6ytVlm9jQrTqq6K1WqSngrXQzfFu+bWneJ27sYJB0lyJZKxqz1AsHbwvvt
gLCnh7Sqes4I69zKupl0snsaeOssvXCtGYH6mKRGeP0jyQpQJF4M9WFvWLDzN8mR
4zinTyTww+bt8f3AWxflhUyOjte6tumRbK7gT4E0Bh2JxvVTJYhvq6E9YMTTC4PH
SymQXlONPn6g//7bqsZzsr4tWIFmZ6LrcvC/3CeprtRBm88bNltTaLwOeGCLdZ9p
gV5ciaBw74hkBfQ/cnHp9cleBeAyXTSxaqcMrf1qpghNBp0yqbrb83gSGiGWWvKK
6uIOn7uHuy1H0bMkDgHAy0Q5wFXB3DZWW8VHfXYgI7KHg69dXL5lzyWU/JRDBPky
05UYnqClUdsMCXc7V6oiGYWDs3ryZrzSghbSbN5MdVXAaQJwyeMC9Flcr+KcA1WH
XKHQxW3EDPWYp1EQ1n8fvcDXmjH4akzR01QyQkxTzRWmJMMYJTu+GhZ/vHJ2taHZ
v0YMnszkTvIjrL7M/I7d9tmxc5xjiDnlz9i5bB+Q0SiNvMmZujW9F2W6Cl/Ra1kM
26NkjALFUiRqwsubiHHmiIiu3xTE4JMlsc+jX1ss71obtia4zv1eObBHKEu2RuSq
A1WzPCVR9Iv3Tql+QIKsjkTWfv70g9Fp5R9gdvhb65tmLzp1m2LumnCK8WJib+D6
yQO9VTe3tyDqFtoWe5+B2oVXt0/WK8HyHC8c+uGRI9Q+1UiEjHnk4ORVZOCRqN0a
OvsjWG7mwHnCjnwCCM5NIBOu+QGekIFKZiEeQ9z+G5UTT3KcCo67tARaHTR5FJp5
Wzj/y8Mh4E3A9mHBYUpYIgLha3P3OFYSfuTggQXwb/W0gqPApz5lCmPZtXWV7dSh
5jhGqbCoZrB9eySM+/gtm4Lb/kPlj364OPLUO5yttJNqyMaDHf6VNnyCWiJIXiMB
uIpKOuSB1vQn7Ame6BKbT/OciPJZYKg9qRRK6IJNiPXO6lpD2IqAj45Z5QlG8ATP
Jt/UlWuifz48JA4IJVM8qnsOBip4FVxkjcQwzOuu66KTYPBmz/dgIc5HlrTRw2sl
lbGnkMPENF9fanIFFWk6zdNjrnXMzP79OUOgccQw9U5SugBPej8ctST+39ef7PA1
19CfvGcFjjTvsrQaRbxnaxJ3w9+kP3GdjKs28t/FzUycMVcHmxfbaqZ2B6gYx4RW
fWfVjPa2CFxYMdO3lcTKjozQd3ruj6/L4xLeh4/2ZRkzsnGUWWFUunLcaOd28alJ
O5yHuGIDqyJzXNzDhdmVvWnk/GBraBtkqcpkbaVymPtedaL8cY1o0hyfxSlNrwY8
8Ke/l9ICnl32gtA3ht+iNIkw+jlJEXsqLoLU3GFJ1urPXwnpgVepZ2ZEjnZQfi7n
jR5G2HYs7Cwzq0KvtUnbyyleVYFIuW6ix0M1Sa1xO5qy4FOFsjmIURTzje/HxNjl
gDprbcoinLypEVYb9npVVs2sMUx7NWzGrxqI3y355kt8/NFA9z0NDT53KBT2mibU
RKontJdbncXL+bTFHJVaqhzoz1hGyPA1oXWiWHi/5mdkwfFPMAyGyprefxwu0jBa
wgPEnkjVYdOfbE8fBXmlMoRhFz0noCzEbT/IhJHuoL2sBR+Q5bqCsvr9WPlApbv2
9HYbuvW7UTgrKlI5ECt8DaQc2fdvgmmYY2eF0tYlp04YEkGirOi3UzqCc0A1cdLo
XIXOQ1ZHyw7z5mE5e4+rPQcoUOhn5Y1IR+FB8ixb76mq5ur8UtQ26+jcXrqKAtz9
jm+KlYfxTe1XG638A6MQiO07lhQ0UzZR29wKzRWaThwQht1ghM73D9wp4IcxGZOS
d6IzsE73yE+q+uc98n0FiQ+mvnzzBRot9BxExfHz3n4K+lWFaO7sDqgPFPQc8Kfa
9vNXM9dfwPWtM/OgMRgH82EdVeFK6iiws6Rw5PNf2FgaqgbWxQtiOQowhG/9DcPq
anQ+XmGRSMjaYuupoE3Z5h37rT7J3g4bHNnpA+G/OaRK/j8ansNo8WGo1HQhPO9p
JN7DDOiM9+IehZRLBwKD0dCDzi8P9wUsQwjqLFz6aRFX3HPYtJX50Njc2Lf8EjoP
jKBbisUpzvTXK/9v+6B7mzX51p632OTvfpJAk6H4nigeVumWljeUVNhndtMYs8i8
Blbh0GEpsjI/54JpTRDNT22S4R/NELT+8L6SVxWqX/eTearu1QO6skEjvrBSSNL8
AQTunBJ+oaRLOApRZX03Uvk83AIR9a7rfAu4K7XN0S5m+p59UZkyJufXypZSveVg
h7WS6aa4Ff7OZaUwlofbUbHn2NTO1iSU7wk097OUjIZZY551R916uguQBbDHxcIj
LgdeiQnIPY77pbtCl0egeBytKPC2QKp6c+P4v2hhHKnwSh3k17Q2HQBW+FamQRQx
EVsatD7fyS8N1GYzwRJZwBdSOG5sMNe8PBExVERJ3k+322xanKEgWgApgEkWiqcK
FDi8q4NmRfs+LfsjKMAKnn2lS7Rf26CUfARiE/b3UFKVMkmlZ1GptSA86hE/Hb6S
4rlLXUCEPEZSKYWs2UifR3UxzY//ls63zBDutR0Aj3ofsIrAt3LKLj/EcXuBdU4J
LYuxEvy+1FcytA0CU03tIDcBcwSBEa7h1kX20bOUAZO0htItIAd8TSl4rvaeH/FS
kSynMyyvg3+8yleD/uRXPVNrcGyD4yksF4sniHDcyWvgOpwam+BiVk68/pBw7Gn5
9p2gnklf1IhJDN3rm5oVEw3O0uOFkYNBe71DZZcioP1gZ/vHn+5xIZbk+M+abvCm
+chHmUzr4VUzVFJj7VrbuH2zfdEhg6M3+H1dEjEMPo50uvlg4t1oMOwZ+PcOZLoR
2JT78f1bDL9jX/PNN875QtQq1TWbEMepgrcRPm3u9zP51JgLXCh8MyUJ5Divj+bt
N3uHlpDJxDPra1qk78FJCGSTxHUf8gtI2rzMbuD7WkBr0I9eaMei1+exfogwOhnr
8ZwekASC93j1DGGFYSrB3HaHJRuNoeVPjcQtCp9/FK/Oml/Xy3Z2lHzW6GmAKCj8
V0IX2xF80tA343mYEiUTou/s5TqH5ToKjJHPE8k2RMNWTEFXgynryl9bmruDraDk
OBj+vOH30mhwkOrkU6Q6OJzadti5P0OdLyZAgkPB9k2X5eGq+suJzaSa2jzqHMYT
AP0kdo2VLQWl/PjeI1z6AwkE7MUmHuwkc502et5EooJ2nlY0/dFMDuLf6wBrPV9U
guMv47NHyaWzRXoMfYm07jh8nt5vO8RA8qCXhsAw2m2Tbr6yqQWajFOTe3zpWA7h
0RVh1p4fEYaXVXZjZd9HG81cpFJVVxIa0hOpI8xeaCI0/YpBPHWVpmZ1eZRMYmPq
oaX54YB7iYni8VvnoG6okHx3zoVGIDvuqiup1m5YkL4IC/RGu4Cr4Kd2It6sDug3
bEkIbIrO5a66+ZVcvMTq6mE0mzrNg0VzreTsK8OgYsaGnbZstpJDEG7ogWwaRc9f
54QNpVBcZn4z0BDBy+bSkcQO9OG6eRqtGm/NUWPYBQFHqKP6ilESzV61bL19OWvT
N7GVmtcPFEbGZzDFHdNY4qRpbh7riyoBshH6lDfb09V6yOOvvZsvFIJltCzKCw2p
5FLL/qYtUpgSWCylhNrPnw5U/BTOSsCVg274fcnfUllty2kHLofUKhTtHqeYIJfT
4uw46Hf/AIxjgG2r6YyXaell+0BASHbLMj4jWy/bQJsML0R9xsUDCbESnZNiM9fY
6OYJQIvGT3VcR6EUigC2xZ+hINnb8x5Nnl+ZpXK5NnSdwIquGkqA1+C9xpZiT96B
1b7g/J9nb+Jk4EiFskmmA0i5iCVPyn+fgWl87U3DCnS+kyA7SztnoojRNXkVuW7c
cLkdXvqU2Q3kdsYcaiMF1pp32WwhTQ5N4XKc6Fjoiw/estgdk34PtopdayGcV7Nn
i4C8eSvFHCAcCVPdfdASDQwcBPHsp6pdP2HbrjD7pOBBKCi5jDi8nIHmVzLuDJbv
uJo96RvnRppvg6fTjkqEbAfwiVF7z9IJLrX2ZVK/ksxxHtgaU7O6oJYM7rpl1jwU
w0L8QpMIkE1vuApT+VhD3c2JUILAW34zp+KPM6XxawFdmP1dS02dWkxd+SiAMt9h
HTIvHRNc3U49ZGh47lIA9ldFs+RSWcK66uj3X1rrord8lIrEWWHpBU/VbKXFrT2D
iJENhivHm2Dw7rCNFf5BKYn/DImM2qLm0y9/9OzPBSWOEqBh1Goplg40je/Ueupv
FvgDbumPaO0Xx2BHxYO1PPn7Vm9oHP1WPAqeuKS2pcJjndZj15/VP8nrXsiEhIxG
MFMC6HH0Rj62geN4wDUQexC548cSjx287RVc93dDKSSAUXhW2nhR+nz59buBkBVE
7nBu3YnBfRfS1iOR1QFP1XJjSu195+j+KkjUCIUMJFHU2u4SiNHRrJaXi1kbA8r1
uS5pxVKD7c2CogwDlNuwr7/vWivR4JrSgqhWbH29ul0Hu5zOM3vZTKfdv6CLqi56
MpNboCXQMc9mFvShKxZNjXJcxnGB1Ttn0Ldi63mOycWr0Z3RRW599nkl3zJFS53L
LD/cc6VXuPhSr4kh8sPb0JlKzEVUCsYXM2tcEPRjPzpdqrkXCDhUXvHRmZaWxelQ
qVpNxOW6OGkyfZ2s2+rHmGfWTqeDrskBsDej8BZRlEe7LyeRpjUI3ZDmRnSjq1nW
xzFSUsqShVo8WLPI4lhcnStr7ka0MGRQZw5ArvzmKzZbTNJDE+92thNKJ4C4GOZu
mKKfK52/uSZrphZpz2exShOukLg9+CiDrcauiKMEDV0OJ3hHtfE4xf3UMuXLnQrz
ttN5EFDHkkoAIH94xEdwUFjH3j9rzhbyuZ+ZFEtPzi1K66rW7ZLvFEStPI5FN/6M
NEJ+sPC2CK+yNLht+od4l4sQAATMC7RVZUr12y/nM4szeVOfh0YzT5ibKUaNIs4e
ePqWsQ7092UQL5YDrZfclhMF8RtrmhkC8sbZ34rlr+8jnnNG9DrGcPHDdiNVnOWj
z12Iy3wJdoVdy+LtHiMQEeR85ERRmaeurR+G1YIZOrSiicHgD2Ye2Jvo2o8cw0S2
wpcmJ0l6Ewiuaqn2REbdjefR47jVRhoq0jpL8cI2UgFgmB7+OL4nZ1soe2xm0ZNb
UZvlLY6I8owsNHMFoGksxC5sghs9LQOtPDG4BwGoKgBT0gwEHpgiilYldV2PQq7i
NRF+BtpjR0AF8Jm/qRiCjQvSC3I7J6F9Trn8PNqKEE8rTAF8wKZ7WHm26ecLbuvQ
w4ePyHnrVzbdUNwMYpqjneVzK9PO/Ydp4fxkjAj6o2D/BDPBgplrL0A7qR278AK6
gpPxLjk88J6723k1l6dlvjezW3kB2HE/+XnteJCIl/KPbWS83bVGEPGIKwAuScYr
/l6WVEbD9rTpLlqw4WQTrufoShNyB7xjmKx151JMJtJuMwEHSt0uBvcFu/cKIU4R
QA5SsAPmjl7YpLGVx7kZf3647FoVmCGQY4zehTWSy2kiBrVD1OeNFrl5lyKFnZTc
SF4mX8QUXIOLcFyHKQ0Uij2gZ6X4wNPSEbu5tR6450IGKBYs3SIcUzO0qiJzgAfq
Njz5UqcR3XTtf2dTzpuvVKhLqTM7gv9eF2bI79ZMDcyBYLOX7fCD3THLKwkP5BuQ
4LOhA8e4M+OztoHnxNZ+Oiv7nW6aRtwPN3LwdJOa47cWk5CsXUDwDFbkePzqlgur
dQ6BJ1WMaFynUl88JBWmJA0r6JLkcu8m4ftH5snjtNCRaJtRqFGaabymXimtLERU
y0VWpUGNzMYFOGdb6VX27idp9q/KMNurGFAhDs+GZiyQxZ4ecM9kQZir/Lcpqdsl
sgHwF9q+LN2PJCmn3muZxaREAxPzbdyQrHKFjsKEIRuWhDw2XI+vS6Ped+SqdjHv
2SmK8a2xSsPuNHfHIf+HfIQMG6Uft9gHIpNzoNUCtm2tpKrpIqt5OK3bvav9/eJ5
QeAWrbWqzQFUaFgnjB0rc0+dnI6sk0l9COZA4jAgxIo8cr6mCDrMzo/430V2dFdq
q8B9LmM0RsU8aMd5OD2tKrEXLgI+5saC1SGbW8MuUPaqcxwaFa2VtP5IEHP8BSwK
cxEkEwe9+/HkvBFx54c2bYzdM/1PyQ2PKL97KGHW5+PO+0GqARYzsdiBvRUS6kw9
VxCVoW6he/82l2D4SNoMifnyebc13CZSITKmmW5Ms+Gv0DPnB0M6tgGkg8W5ONtQ
G41kiknmATYtTrH5AB5zwHnFOLcHz1ejnOf2OXZaSzrOZzhyXcSBCbbpHDwXOGrr
KfIOruJ2085CPZJjzxmFQyqxUVAz8jwV+fVr8jva/w+D2Ye/+N0wGefxaa/yTgyf
rSPzPVz4w1SseKkmCxrbjmQqiZfztBzuVu/CK9pe1GRKHtO7M6Y/tJB3XP5qhlJW
eLvQekSk+1JE3Mmw3xPXI7TtFD51FrQ0QKLZYO0MTXrfCNpkBtO2w8a5ZomZXPv8
PO1kGzXb+gbadoG2h0FxZFMGo3qrbTgj9ZEoC1yy+LBYYue7/w6/Uj7gigiF4nwH
YhE2mM+EZjVV/FHbgrQ5bkmPATQfXLo2HYT/kp30oZdebm8FDlmj5sJE7Ik7+YSZ
8JBwf+Yt9NC4CjliObmCpL+qJMs1/MaPhO5nl/uUkltBbaulqegC7n+wq3rSwU15
C3DJjgByyqsK4+tEfqeE/ABwP/sbN/EIWcPnYKIPs4i027gTSVpUQ6JCJ6xg/z3o
zgFcBeUtG7HTvgyAURebb743uHfZXysacc+v4PJfJPWSDI0y/wv1YD7Apg+RJPpe
F8L5MHrpDAO5bxJmp+dpgmW3MAeRmU4ZrAfnVeaCGYW92T5hO5tm5jfMI8gh+j9U
TkUadN5m3E/MJ8dGLI3vF94DRbQUmKXe/wwjNoBrb8QbJiWaY5NqLVvD6yuMagm2
TyFmku5i7ZaZoX+rLCrvvTsXsDLamCbmGogSdI7cRwVFZnX77RHpCuY/a4DqbV4m
BYI71/46VWCaIpUww2DHkP19j6Suki4+KV7goIdDXNDPg7Od/cOQfOH3bLJrVpHY
lxZAH2DCSAwDE2swzq8RZqbV81XmwfaRH3o+OLCNr3vADYlL35rsjchYBqpTkoKQ
8sGoucLL9i8/FFJJrQI9UsRgmxctY6tAsIS72T9lilIZs1PJPChsMWBO8gy9NDz9
tLYOHp86zgc45Pj+WGH1/M5z77QDqsjaiGW8kvZTjJQ7HGidS/KO2nSlmnofBzFr
xfQJrxP4/P/HdnBmyMeFB/Nkvt25nxp5ed/AxyHVR3bZNa/XkTw9wHEqmpqLqSPv
aNW4KkVC/IV6AMVHYAaH90ORK9oPm6wev/M6yB7kvpVbo745V2zUgjOaePJg8o3D
4fvUO3CTgoptCSLTWUw8NVSVA5iJaAWSMhtYpHNnhDGjmABWpyNhDi8aZIP7LTXI
N5UJ/1YFXXvPbf0EpFlQZ72BIvY3ExVpMuzjH6+cwXnNkOu9Xy5JgXQKUBakPaRi
RdRMCMHK0trXRb/4ubx7RrA+UYb/OBMYdnZuhB5sNstrWc8K+7VqxyRAKAI8XApL
8prpkMt067yUXDhUHSlvgPM401KS3GoKG3z07KjWh2fSYRHoXT4GTLoWQ+ZkHPoh
DAnPx+U+/CNp5nNDHlODw4FsZW7gWF22lX5a0C9t5naDlByfBLCewS4+hZhqi3jh
4rjz8j8dUN9ftrTMKGshe+JPN+aSMcei19OHnSWKa0MeTi2MgK/kdolAzN+jqDIC
osH8/VK+MtozG+eZeoeNCIdtS6uh0JLZxQ1xG8ydOvDmoaY6Rb9nHhl+gQ5hEJGE
6E4MTzpYE7QtaAyaaBoIFxYat4ar16k9uUCQPfmvxowuUNTnMciH4BMBHhpW+jsp
DapVyGAaouGzaqpPxPT97rMh6asihL0nx3dI/bK51I9cOWhsRcKhtuggFVmlFC3v
fwLC3vcX8D8ZnktRE/edIE/4v6nd6jzE3kfjQnXAZRN87CLMx5JGiH0oYiGzQC4B
9BrEgFUiirrLd0e65qAwdQqj7EBQYEF/7c1VlX5OTW0X0CoXY70par7NhaR9YqYo
xPkcQKuVo+Z6yMhrffKkAXICQjWKvRLfGqLY97HXr1FvBqyUgVTK8NDRyKN7ktsq
1HqazTXkAAuPBHVrBAYXDpgGQyp8tna91ic1JsCKro38+l8L1MHOPvhoBvxE9BFG
hLPbynK4nfGL2g6Wru5iDk/nkTxrPlac+HFr8EdjA1N8KHphXxZ4RhB999iNCxF0
OqdhScdwX1jxTKBbpq84wPeGH+Te0NrHU4S77eDMR2FgLsrqUfT8JtuT3FViz6BA
4Pc9oooSFhq7TwAlY9RNGHd6Yul9KuwzEiPoSTRvdKXq4Xo3DiCR6PFaSJD7w+Ud
7KWw4hfDydl7JhRh9ymx9zzv1Ri++YS5Y9aUNv7vGoEBStv3iva/RUc3+6+IKMF/
Hc/4svDxIbLEooGyoqq4FOwJn44N3/a1+/1RrTwSP2xr7wM97bKCTIz0qGRUir62
6sfXc1zagauh4IMKik8FxfKWrY64c/1yDgY3T3M26yoggnM3pArRT6VfZVBFzAbF
jyAaafn6cM+/TdioMti4bOvyqeSh5i1m9y7d3O9rudv10JWKUpwVw14PoCC9Oj6x
EUtDYH/Yehjt8ccdoUblkf9OnGi4sFe21P0wwEXPKZT4b2SdoPztbRPhJxYAhjMZ
R4gKTcczUzDkXd+OhKNVVzCLipoJjLvyztJEJFNA2QVnkuSSt9VGmbbu1RTIFmjr
rslbyPXnL2Z+ouucHGDBNE3kKxmqBWrZu02b8rMnB9DIoasRvHHJGuMBo4Qn3+cb
UPqw9g+SWekwYxYWPwb1+WcxKDCP+Nk7wFTnD5kU7rqDYnTzDDEhLlTxnS67yVIg
1/RuSP7uTmBbzL1pGW3/AyMhAmn4LJnVRI943mZm4j+gbWV0T0TwaJJZ1DnF75yk
w3QQTWuzI2lFRBWdE9B0T0622sQeMK4iEQNKLWMPMhzt5qIc/WO1WyoQEmtN6ZJ5
+XujNGBxqTUJTtzSmUkQO35pAIK19cp3Ym2TzGXlfJwVUsA0ORFTotaBAQS2uER7
DDE1Ryatatn4dm/CRT0agV3cyeCaPAsPFIUUHZ2htKukw9SoEup368tSXQBV4wmH
i1BtwFD/15bC0SlvxHuB3rwVGWvfnG+sziIzc0rw0PZU3VON+9nf607kMQ9d4efW
9DFDbDoXZkL3rUlNEa5tq8VvlFoFt4JkwRSxXxK+dGoxAI4DlS16iWzlfLXc+nZO
uoWiCVkHf7yoSa0wKG/E3qHNU7M4KWWIIn4mqW2K3cq/akKvfSClfzCqylTjtJ5W
NOvs95HLXGPV+YOoJpSW7UX4UfdtyazQNYBAsgdNucOdtnlsBsQ0bx1aVLN+30Ji
JdgL57wVPU9I4MPCQoYP9ybcu6HMeigwN4SOaK5ekDzTLg/jYpFw0z5GewgNgTSe
3dZrDN//iJ/PuG0QKZNwTN+uK4z1EycqOp/sV+EMn2Eg9MmHvRoW5aez71wpf44N
yJdqbLJfKvbjXfCWPgRM+y97T8D1PP71lxyPYVL5NHZ9dPvEUE9d+jDMW/EpkvRP
Q1bkhx1CdxrekYGxY3BXwiww6rZCvwWz8EZUjM+kHLfaBKzmWWYZcx1/sNwjiUNj
/Qv5ouNF/CsdQMwS5KR1mXlhQWCSstcvGbXcqjFVR9ceX2fE3/t7HacwAPe7tjIc
efoYsshAofInJI6PsHySCxIMA+CKAEohg8wdVk+2ycsv+4zGLqXNsiSEKnwKPhB5
oaIPoXBUf8IhBoRrX7vsoe0sHujQKfs1ekYeATksceKI9ljgqLsqRYPlscqOs9y5
pIIcfdV7NFfu8fZJS4O/Bq4BGTjgwGgfPRblsirjJKdFEANwTA78EDbwfHyRtXco
cEKUR5pWOb5vCYKOQbWpwuaNED404BreNR2ma0F58wnE2oRlmEnulPHB5dbbrH1v
LngaUdCaE1t8/UZT7gWSqGsu/L0+9GTSQIpEvLxpf1W0jAXjtA5Gphh5tCSLJeLP
amwjfS7ne1MOdhsm6q0Kt8O7QcQmpSvivaC5rEKqRp2GQ+z9FeA/MPe4+jwh9QVM
wAoW8D5v+NsEWGJSx3l1T99fwHZS3LEZDa06YiC0gtcGbP+DmmnEZ2YVvekh+mNT
PcRrI7S5I+AoOGyVKo6Ni3uS+1kVAVupzou7Bq4VbdVxA7SBKYZtcDo7uakn4I/d
SAmpgPQtWvHpVEVyIQc0GCHbOkU8qVP7qLgM0ySzWriq/QzxcCRCPxBAJmYldVK9
26Jk/NZIXNmrCbt2kKNWlcNLiD92RAxjLttqjXlKjknNBdYon3SkUWdGYHLBfD21
WQkuhl6BMaDMwSoxF1BiZzOay+sPTP+43QAwAUyhvmy4y4kiOuAzK8DGM8J1bc3V
28z6ESAtg+8CKy6aY1hW6eK4ctmwr8zMDZAw5LTJgIgdyZGVRP6TlzPSpU//9WBM
IzQ5sU93hPzMX5sxlIFSV0steT1iTonhEU1H08MckRVMlu8kkOk3jvJqS7y5efCy
jzcv54rv0LmhJxmu6dI2hsrmCMazl9hrlzDV93seWWP3Jm15NRQ+b/A9UB80wFv9
RUWvnWW3IrEAtbZFmJuvqM1qVuH6GjymlSpOeBHmadTs0MmNu7Nswg30WEUvZ+J1
+YZwMlK7sEEin/vYjWUA8SEv271VAhLFzer5g8JhsriXqrBOnI3Gp0RVXdjkSe/B
pkpI+ldAr/qBNyL3pDk8Mm923Y1IvrLW9TSqorv9S+D3gOx8wLXY3uP0aIhZ5UiV
6j7MA8wCLBvSOyt8PavnhRkIalx9gqDo1YOQQZ5CZFa/VvUWzOSiErT6mGQ7pBcl
REf9/TwUj1eGDqYDfd3/vMvo5pZvbBR2sSTM8OmFJd8g9YVPNbr5NmxScYTCKh1C
UW2VOfO1FTtoIZKDhmVEpARzKA237XXismhws/UyvunsLD+KlM8DtFa4Wu45P1MR
eLquZCyRT3KhHonNogqgZ0hUoziAA9adw4UMs+YS2xbvkwdqXc9ETWhLQtTXCm4y
1Q4MeCbZ5Adm1RnybjqSg4pDYdSMU8hclp+Zrzs2ny924M+3ceb3vqqfx/IeITa9
ScJ2FS3VGiyQVaYsoJX1dHjBvhzV+ZiRHXtpOxey+awKYIKCEZPtfn95sIFw/3oB
ofSmAsTq3golVUXZFrUAugSH+6O0+fHTnLTUO/Cp/5uwO3uVr3qxWVX672qscFvq
0lJ3vy5BU2ODAAfRuwNs7CK/It3sm8X5AC2o+BsTkAuLsXWfRsLSayJmlYbo50vk
4VzOF0DdTTQ6/rcxslDyAJqUucpHNWp9N/7GCbidjLx9qps9XTPENf3ktrVuYLyT
GbawFLXVaD8wuQkx1m2WbczwJ6FdFQtYLlGHLkGOHDFuyC7UGn03/Oc3hFD2U5EK
9CwvAVBNwkqao+Kssisv4Tr739YO4ePUuVHRqhdGGBmsYq3h042oqiyQqJWRo8ye
/Zx5qA0+l0WL3XODSdTHajVVrTSSoslpZIgX5stxGpq7W368BJ7+fp0bjQz+F8Zz
p6o2ZBGKaj2sd8U9VvDHc4EYAEohOFN5EobvbtJF5fnIHPLNpeYa5OoOTyZhQdRk
oxhqqVb02cdN2FbY8Qz0rblRufmFyz1I1a8J7gMJ0wu2pwjZN6G1gIicwWaJUG/A
pH2DigYbpRlhAPGDbDVvXTen1ep+GKUNDwYj2atf93IUmwD3BdIurcaUE0nTUbZs
So8DHxpkTmdLhmhemq7o781f8SPpp2+oPSOnXnS7fFzRE/HfRhsTYB5pksAFtafv
VQqG1+SB/8IMQPeVwOIwoqjkp/5SaEnFAARsrqBR7jFQsGG4eVSdtIIxSsYcd7lF
oAb2TugvKOOqOlGgKLHxQAVSwx+hoMzD4zEQ9jR0FhHZMU8lIPeU0InRe5IDtHuN
D/FmWUBOirLTRq1BhvcEeE4aTbhPUtduEWWwNOV41bsVEWz9Lr0mg0g/UjrHaMi+
Yaf9Q9mSGKR4vzO2ZbifP0E748tmsOOulkH5PpMMW+3qemRCo82Ifd+E+/vHlsy2
Co2fwACDRw3qvlEleP6rnEqvfOenU6HMt91L5kY5NHyVW6NJTTCHJlTjf2K4pOlD
xkQGJwafQ5hyzWh4nBOBjhP2x+3waeIdrA9mtC8u7zbY59q8u6ektEDB9tiM1NCI
xN1KpxizIE3QGrP8vcyfDKWbKqEGfEjmDzj2ItIAahZvaiaCGEP86FADIS2pOvN4
gaoCUcJZzUcmNrmPDUYTVQuzSGVh0Ft8SArjZSI6PdzO08zKUxhSS8OBvp17luwC
+ry4diOayMnLVUwCj/yqd7lP9q38ZP/qbkcx7INJVhWPx6cAZKh+JVfycbiB7Rak
SZE2huAlqT7n7LCyAUTyRNaE2HyM9t0Inh4nCQCy72aC/nqvDovmZ1173+suPtDQ
/GGI35Reqv+bmQinxEBnGCiQ45NFbgCOidx/zuuHxWkzI+1LQqAJRXcQEkS0Xta/
Ma5oKn+MCL4fw5QsVRoWmmUyTwdOaSuyxIsCzBmXggehFRIs/qsbsFT3RHashyop
zoEerWaDmvwh1eDGstRXm2vBQ5MxLMWruVi0XCQwhW87sKTDugppj0A/F0gZzppn
+EYj843cENxUVtdnd4RXJ/T3sQydiGHdL7b/lO5bbYmnfajTn+dbGfc7Yf8XYtov
bUTMC/k96mHA9kkYSPFKsEdTrXk4jddVaaUhsXomzkjbRZlNst7f3ug6CGNZDW/K
tsintTtwGptZ1ORC1MIu/9ZbFrNueuNmVcCmIcImTUEYgt/+zgt8j24Yc16A9ghD
L8Frb4Z9fn2PzkfWOUxWtjZz1i4RemgoJXrsvB6FUwIecqlM0d2E51jateK4fB0x
hlWt+Lg1ldwZm7nWJB6ScfWutVSYFa2MPlgL0GbELv8iVnTmfS9zI8YuE/+TXGNS
xpTdFKQXN+/NFLdNFlJoX11uZ0fA4lKXmbDWh25sJiD/2yZP63qpWKj7Eq7PRNcq
8Xf6OFkKvl35vZN0W2+ZFYvJU1+85yS9/Nx2ZQMuySTPLd9QCFYKsaxrkahn460q
jkf1SaH4pEdyItdsWDMO8RLJF3v7IXEM13G9tgPOqB1TAcxynAYlZsOvJh2NlTfT
cEwsHFmyvixKcvqRgT4MN4BNvWeosSVDertSANj+G+1BFQDL0TjSfYReK1CFQLeJ
3rz5gTXmkFT4GAGcO3YeQy3n8BEAORLa9QrfoJTYsC6OemD9qFavONRKORe7aCWK
ghOm10X2jNJIHf3v1Mgr9+PuxWNn0wolN3peseoVMBl5V8qMDtFwFslsv5plhfhJ
xKDXOb1g6THaW+M+YsiaSngX4PtcOvxx98NNxLvV63589qXAWfK9qEFVGLcU6XAi
EgjXE4zErT+hnxLVk4zIJ4d9d2FdZSXFOXTjdjPBxLbvkYxzmydC0rkDh1J5z6+A
MfVt9peTdC+4GFfg7ab8dkLw7k65PKIXtjlFq2FFezNXwQknIvcQj4iCPLMZMCG3
c40G+fv/j2jsrNEZk7mLgtVnqHYjPPrtvgQ+F41ARXtZC7xuBGPavuSrOYXtLu2D
0ZxWtfUa0upOCaHgnKHtu9fFJUIUOnJYCJUChnzjZs5SMNObl61H9bQa4UPeQ4GI
ptd9/S+jXNO5bVvUgbmXoeSyOC4GNaisLJnY3Pnoheq77hGXv0Kg0i2Z/z5CJEnE
bFw5yeheYoN0eTy5ubKtalcmuyhNfo2lUMXZz3dQRRozxilwi3fWsoMKskLP6ofx
57wqgV8ggoR8UsA3OgRfIWlT1cdRNdRCMmsLivvnFJsndvI/QsNP0l1DfZTYQcWC
u96Ktuo/0ZY3PHjjhztRm67xfLMYzoSLyg/qq2goGtrZp1KAy8yq3JT+nOm4hdXT
pbXjMrc9U5Ts+LsBCvzTFxemfjNKTKl7YrZUgwAGXGcIz6rc4uEIVT6MYnmwuno0
MDYAB/Pk4490z9S/uuKvUSNi9aMmEuNoR3iIHsU6J+ysTZTGYJRODQblor5jkgEh
OduyQkl3Ok1BxrAARRqXvMUpqKW53dKc/1GGnmP2+YAy/Kk9+2/on2Esj83rqZxz
WllArahEDL+sT5yFpvuDoNGtArxYS0j+Myb+ri/GX3sTT6ikOIQzldK+IO8MpkCo
Eb3Czzcctc1BOdfcvgSlRPc5uvT9yHR4QDhaC7gMUEP4oah2QMnhza2dEDG2/ljh
40+uAa5A6YHHEeaAm7QeD7t7/VR6Topb38n/yv1gmjQ1WlKheH1Qo6pSbZ96Lt2j
G26NBcdHQGQpK+EQgWeW2gRonjo+gPuffn9N3szNO/fEdfZPhqtTl89Ax7MAeSzQ
5/7Ka/ABeOh/7sFxIu9OUeCcbaS18RaeztoJfth8Z6Xep293VtYB77NEwfh4ebyN
Dzd/O6kXXYsjPSOooY4nGvp9qheqSrUAzC0ohjLxzX7+ZOGqt0pBnSXobr4NH7PE
SITGvKnPN2uTcL8iFn8Iv/rVM2Bh8sFF52rY0InkYmDwu5SvyhkTxhCN5GkAgtkC
ofVaI2LXPNmWqc5udo7eJtnEI3rQteYKCuEFly/xOCAZMKyWm1/ISRMAyfopr6GW
3PAJq1G2oUNNIPZOo2wDQaMCaqcFE4owyQ8LNrZsYK502IgE5wjvDgyh3YTZaRQW
cB/QrqHzETyA5p3wMuhuR2rYXRyUhxt76+al8h6X3VbKaOn49jRP6yeYtnn4Tsoi
4RAH/dr9CAuFhegTuNIYGnFefkBoE3UVutiNiA01wev07nuzdtWGChJIxlcPA9Hi
rQvPJ1hFGgZ7FlZi6NXcEZ6lIpAKjkBqq96WymwEzJo7js++PLrIjHFZ9m7PpAfn
YXJvfTQt7uyj6fhq5bD17YDi7woxArCXsVrBILATtOWHghyu6FLHWCuLEX7H9YAt
d9jSFVSKHZsXJIShYl9WzBD+aqi4SfTkNXcAj5+ks2vyjJGU41y7MnNM0CHUj6Zy
GLA/Svsh2sQRoMw7jtFxsKrkv7E3ps7mwhd/+L13XL5GPzftBpRMfsIntQcMtIua
2ffa2/iiaapoy1ZTMYihNEoWbp77xGCRu6N3FBDloG8XAmMaSJQTHxAqUayntkoY
2t60bKnqjeerRjTrz2idzfo7wgiNNQByg49vQteZlYpWFrA78CPR/DVyT1UhU8H4
dkC1NbW1qKojklqMVQUXjJ7K+YX9l5GgeUw0Fn1mg0IruCSxlhz2MgRXkM7X4vTO
HCU6MyJmNT8ks92F7Q9s2vrKcPdi9k4vecnBvKtpLTM+5MwMqPhAcujZ7eY+oaUg
KXvdwB3R/N8l0LhtSSUDm9jUFSBiEhv5UPndp3kKLvfHjWoect0mITjE5YyBYyCl
grpRU74xHqcFsCym3QCO1tQJY1D7DmEybqBy2IHHqmMxitNY501Iskr+qrTU7YD8
E4mOzKCvYDAReQOCGOJonl8y+ACjPARS7ZSw6Psi3zdxZAT45tburek9OG2jru54
Ldr/5ky1t9+Qh2UbjXChiwrFcmavyQgWQv6ocTbaC/wm+70S5AFlE+sfxFdnvLnp
e5z5kCT/FLbpu3+zJjEEqe2PdO0MJAe/jOndJvAFIQLzs3wuY8heK7Fb7UGZMrNX
mwEVi39/v2/80jMi4cxbbELiFv7vRLYxy5LWxtQaEKNOslhsuW/3uJucmjbOuWXt
i+cBuAbR852q17Pp5716DbiraoOz6INDpcsiAbUx70WQ+E7wIyi0yUH5MUrrfg+F
cNWUUgKfP0UwqoyRQtKYBzgCwvvJQdKZa9zzmIyn9HD8C9aNOWlW9LlFGd30UUdd
yfgCx21iwUVHe62yILg7jxeO793izv9oxLViMsAoPsHqrWPreE/KqCmGySdKL7hH
aon3VDymVD07SaHxjZaZIRfiYxPir+y8ASmWW9xfw9mj8dCx4fqJg3zSw4yRhYA4
dmpOcDinEWKt+RN61IXPAzt0bQ1X+kvr9sbTw+zooxo25aRCazbpzhCcIe5/iZvw
hXnEe5C9AHk9SHdUy856FtYoCf0mFcwiUcQpdzg7871S9kelXU0HVDdZJ6KZJVDv
p/zTLAhCEd0IHvP6HAwyd0CWbXgNLxt13ZclhNE/ZpS656Zh+XFeKz2qN6wlJFtQ
gt3VXO9r3VLD7N0/+6+n6QtPB5MCL6dDeSxUlWxDDWHI2N21iFevWyBNF6ECmK2X
SY7YaX9VP7yyNFtNS2QAovnp7fHjI9WtxJPggTrOJbW2I3rpIvQ8SnX9+BVt2lMm
Urd78ns/RHRMYun+qsIht6egWUSqlMoPwyxqtGVnCtD0bFsu8srQAd6KIZExlyG/
0K6fuoAaBT42rLsN8QwYFjf6fN564OqioUdCSLmGBH/gmfTkr5FVsWo4wCtV2Kr+
82T0IUduocbO6G7dULoISqVPg3sLw9ag/ltLCb/hu4elJVuRDNuyHMG4jBteK2gU
T8A4jj6B3+r9I11rzXiqB7tzIINJ2i1zl82vkxV6oV6LGB7HXMhNCkT/C1TNjB2h
y5oOmT6QoJ0W0HjlaOylvQnGLYyGpMQ/36+1JOVaDfEZEQ2QzctWAT8+KMfT1BD1
uFVbsV/dgfHzu2Bgn+VEbXUmKoUwwhU2/hYe0+FOBIrg9SY8u++B2TYbuwerhnmt
1WhwU/q3NWkuzlqgb4AKcQICrIJOGQVnqvnFxdkAzrT45ITmtGE//eWvoG3/iMLV
DoPps14YlAeGfiIyDUXylyTfsAniq3VQEJSLWJIrRlHW2PC55mz2n3mzw9oqPVtv
cnIuahTYrBBHEoVD5QvBuIkBeAc2E6RueD5mzSXS7HJ2RYlNKPZNPVjpw3YdCy2o
Xn/MlGDt7jglEomRCVcWW1NAy/X9yq4vOyVAMZNtYzhzjAV2NFuSkU7IMFcSDq/V
7G0ZQ4pHlkCPpuC1oxa0N743+tDyaz9bjdu0KiPI2rI9PbJTt0TOawECPWUPO9Yp
BhlMlobuvFkJpmcfQ2jNr7Hkev8nfeN8Wy04BV0Pd/hNBioA0lyVpbnJa3Do/gvR
4Lzt8cnBl/JYgpcKmR4NXDck5uHBt0arfUBfs/txPULb6dt2uHAHjVCKLkybDTMt
vu+RG4JY0eCl82f4TPLz0I8RoVhfjhamGZl2YzcUQ3eNQNYDnUGvBRi2QZTm9UOB
hUQsFrDiZrOLdsXUSS0wg6nwr5xATKJD61SzciImorjI2Jy+WNLsRfqPwKERx9/P
SBWSPalvBumU1r/17Rgu9bB6SvueuH2adEADhj7XoKyVwYs4PTR46WNJFR/2bUCr
z7pBDh3AvDe3cLQZsB9hgBySNcAUzJqT98ChtjpsZAsYixT/3gHLn/vZ2UXKY12A
cv9k5mbMbicwkcXQ9zBLfLqB7t50So+/uRSNudPtb/7rIl+dBwqpL8erfrle7VlA
OvL40FgwL5FPDt+gTXx/ssFEdhLq0i/PQ5AXD8/xJ0nAa9zkQaI/Ai3OFW0zdJQ6
kaYbxbHNUbCyUgJApKCLScZ3YLn8o8PJ+bS0F6m7Rpfbqs3wLDkqkwtwi92bJTgy
0zkTOq+oZtNF06ZsIJZe0zZaAyPKjv6Ry8orMcRHMwzv1qGTQvYzJdVCDoEvizOh
SLVX47ysSsYn2x1NhtEifyfu+vv1MHyMN4LlYFQCF4H5GiUUc9QfmUH0FThywaHV
tqrWZ0bbc6qsJvQcF+j0qODvBzPGLO8o3yZrVCSYsIfmELcpjYEKoy9E3h/Ng7AE
p2zymd8vTOhO7yFYjfAFMz84wMEmF/kMh/3DVApR52GHgDDRuq4V522mgm3Y14LE
XpRVH5HU+JiU4qwLr5OLn0oZXLsAknrOcYEnjaCdK8CW67NaxOZ+/yxi4YMK8b/O
iL0axewoxwfJTcu/zVT+xfAki13bA4F1TcxTwDC3yRMi7+xsYFNTD7n5P2IA5A3x
nKkz8xf9icn+6W2542+ZjAwvB5MRbNl6vxr4I5UjKt556xZyq4c7PcPgPKq8algV
yzf+Zj2g9rbtu2htBqATFXVDOeB/MCt2wAVkxGO7HEo9eCjs5zSXvjOb5Uo5GYlg
Sspu9z4zZj0L+B8OldqQJsG+M/awhU1yDY7SD172v2eiBVsHKXpQ6iMNlZ2PXVAm
WIGyTVfKTq88cIpxu6yZDR70NrXL2yqHtmBXvQVwliMMZDwcRD823Gs/F7hIQ8Oh
AyfI3w2CWpcoLp5OW2LdXuk+DjnDuHyjWhNI8HkRlq32ZTxPUzexzGiW+gJ634OJ
cndKERPujynkoeI3SSm4yEUGCI774SfLrFRBoOw0xb7Sy6fzPTiIopl+wluMoVYo
PPvYnlP8bCfrzn2xOQG0yP/YRGx/9tWA3jgjzyIpek6WvKjyoC75aOEm0pKQXat+
Cnz8dHkPdmnx68oj9s0MX8UI9dkBMYvB2b5ITHn0EvSHIK7msBVEH4L5+GrQP4EJ
cD6BMmfa7C33ZCdYFnoV3EzpgB4BfOL6ReBd03z+iI32wkfn5JZu8wEBuceFloBJ
g7AOgj9HDOMfE4O8k0Xe87awWil2Q77kEM+m2QQzJpwumyl61l35XcktqV0ySJT4
BDUTd2n2PZUDCfUpGHSnXg7gq0K80NNE1HN0KEti1FGYcDKDmG+5o3n/xIrcvMFp
8QeOSVCd3LNR6lNErNJGsWGDZOvyA6mrsA4mtrdOwUA2iwkxwBmDUBI6cN3nKpH2
bH74aPn9WYrlzKVVGnbXeX3SyiqmVQKoj3XwSnj+1sSP8JIXS9ULjZ/RaTJV/Ugn
cceRRww/FJCKp5zIRxfGuy9gotiBzpnVtlrn61LIhfmbtqCSfbM7+CBo+L+hoDtj
GrDXNuzicSDzRWZdzivSQj2T4q9PuO+xlAl3nbBSN3FJkDnJGwmG0tR6iM4K9spl
30j3m1e2Murhqv7767dT4B0MAtOKw06AXEIRERt0JTekPc/TPY0eiiWeuyUzjnUr
9MAIZPofAxn1n9REM8VTi2xwnZ6mKy1Fs0Fe7wekqKi4QuOc4GX5SxVYUhreczHT
kFC2MblI1ukqcrQ4uT+rJi90m88vsL1ZamS/8CAaywXVkLH1YuYdhG0xK1LUtMjk
M1mownmsXbgb5BYvDrcyuasxawWwot/KxuABHS3RYS+LNWhY98Ra7iYXvpJnTOru
rJ5lfWHfJ/6Gwpq/hfieuQsUD5nSRAPpsGzLTo8Hu3gcnHoIQd0GGj7K3BJfiepM
HJrO1SSdqpAHHIxHTtcAAS2hjifr3ouqMI7Fwipt0GwJynhIjeQKZkXk8JOzxrHG
PXNivH8Woas548WhaFO+18t6IR55NOcGS/FNcM2cMNnLmVT3lpGjJn6V9NNhbesJ
1VuHZXrcjc8kMbSJQa3JfltueKASeEbUvKOHXvM6X6F/P9w9EQSLatiP7YOkuwfH
edtF8sw9uWC0e2B31Q/ZaYpCdtWFtPZopnTY/q1pafaue4OxWk8ql70wiUKQ+UMX
x5bpFxVayPAHuwcpu6wV4MYvqMcv1yTMFg9ojLnqelb5UAwNr1k1yfcbCJLvsMCc
p3WhsFxgI0r93G5VD63yTCUDibORO8tMLV/cYmC8eevRE83a6iUt7crou/lGlbLh
/b+Wh7w98rrsD8DLKOWV0Sb4QCPbNUwu3VlRAgt7O2njGLSevULdyvSHPqhZqA76
jHvkDeaTRpwpVUSv3Hui6soTIdLsqvkALwddE4pylmj//kfgOn8QOLivrfr5EpDZ
NdPJmumjLVjiKzmfEWgOp9CVsvKwoD8VKqgM5XgS1V6W+ABMmglh/nRRmW1P6NVM
e5Tt5hZjqWxYzNDBhKgpyItyuRDJuQXYqr0PGwjEs9lz+Yns3B0yssAxLvUFf2e4
++Cy3VHV47W0bXJGE3Re8J3s6Lg5sjm53Cct/gLJyh/hUitKzDxhvUzi7COuqOfy
Osf/blXKrKQaELh9tzGNt+vrGE2hl6CvRF9wsL5qdaHcZ4TDfVTQ7++xD5e47pvq
x0mGvGZDbDTWEbz0zdXIgK4unAyE3xIUIjjyD7IP/fTQAT0IM8xllvbg9e0XHny6
dJKSdu29Jo3tYuV69dBOSohxmfOj6/ycUAMqGwG8uRMeMHFxAHovjh1gx8t7X079
C+zZkyc4x9pnLBSEQq5h5IZCBTtKlLdLYO/90WTG+OvlILjBcMUcf1VpijTJvBSm
5VzbuxiZL8kQJJEvLfgBs7U+Q6biAy7BM+noP6HEgHbAT8o1xQde/v35nD9fLDqz
y3Nw7xAsiCnjWS5ENg9YKxZxQ80/ZxjwSIEPYeaoa/gEf8LMETT8IcUwPv5IyQZJ
KjNmAukSFeh5XSfnVq/fzl9bzCzJoDit4x0CN1niXO7zSgIdh0sr2fozX9bpHOP0
ArwRepCxEYI5yQjqzLhgeRFi1HNV8k8nlposcgHqOLrDERm3FvrUNRclAexceL71
51SLz6SOgyRsaIMOo1io6SyvZ+z+oZXSduNOz0QHTGfdpwfwSofhu7pq+7iD4U9X
55EvFt4/CpfYWwkL93dT+szd8hAHGjpA/DjsI3P5Klh2RxN0NouFz0O/Kll75D6H
GbXA0FoNyorPU/n+HigiwMp7ar8suuI6qfxLtxbpXkS1N6xf5fL4HK0jb/IMnqYh
E9X9PkCLefVDFq72UFgOiwvALSvEUL8bZwP9S7N2zXvsB9ghn1/L2J1JhoOPglbV
/IRYIrPHR9hBFKDFXuxxiMjO83GMhqq0bNFxBQP2JH6T8eySgPFpmr89QwPWSZPG
s+fx6G40fMwjoA19H3BtSAJ2eiZLNfR2B07PsQvFIhKkZ7qCzGrBBMzDKEYTXPx8
xCJl+2ZIT3HJsvkxhkGOvoR/WslaNY/kDFaAYE9W1xc8+OwnyoZynzoo7bcV1eAy
fohJLYdjwXmVBsNHfYmcKqLG/Lb6e34ka4A2g8AP4W69FhmoclEot++9hBPE4rNN
SIGNF5VOzBA84lUmawHc6Ley3UXDJp5X0g/q/iB2SdTAzJjpAxBHqR9HWiW2E96a
GW/Yoz+KISeNEdRkBX+7eXzVwUVvZ8g4U+NheCGPcOTN9kD9C6ZR3+D1EEouxH+B
VWkWBSSRQKDxz/lRjay8vjSpKJuwS9N4iefiWT4io5VlkjimAi5Pel9qvnxYKxkq
j2nPZxGiqIorL4IJ7V9wv04trrizGfTzVuPzhcnJPMWO5Oo6ztGvRmviJ1lMewlN
UD1nfLU+u+QWYn9StRIGsMNfdE6hJUJZlXi59f8WNitCs01d6PY7lcF9k1Zd9IQI
nTNWaUCsaGhME/GR7/z3o/j9cVVXKkJflUTL/YaDV84x03YDceImAc+ZZkr3FQaR
yU5JrttkPnFsBVFYofgNsec8g5KmCWmtYF5M2YVTleT+Jiyc6Qt0yyNI800fcoYc
+y6moLUf/CiEf3Z6WKAd67REl2R7TCe/wF9y5RUOHnJS3OTY6IBYSTd2dbldTeyi
uW1PZ31WkgWwhOTgePFWctLBWkNVkiom2wVbJjmTZVbwG11LF4wO/jsMwRC3pmk6
qUmOrzTTVOo3+XiyiEqPKNmZ5up/EsoOECIsf9c9IvmJI878xA7N1i+j8jdUbANV
c7/nlAq+2yJVj5bBZZBmng457OBg8giGguSMp2lJca6FCDll2o23UGyXsVK9c7Bw
MguhwytxByUuHvBw0t3cmStEqwuxN4C9tpouXGhZnpNwSjsfvpklHl0ZnY1bBx4q
V35oacd5h5bJlNN5fALh7h20RajPfT0ng8YjCAnDJjbokn+5wT0+20Q0Y9nYH4NT
+o7nb4MSSVt9pM839DfHMc/HK356GOa6Lfw8VgIl2J4J119XEX7dEwDQgEZ50ytW
CxJcyPhmR8lUF/ulzg97E5z4kVWAE5D/haIrzjvGFeRY6lFfIfG5/beopFm3kYfQ
cutIcT5q1/+xeuQaLxJonb7glcC8/m4l4Z18oLi3NcWCj/BhEQcw5IGFtN4bS8jR
wNnwIvFb1UHvTPzYOPTcAlW06o1xJTK9dLXv+/3IUm+0Gei7gbKam8oKEGiw+OuU
z42Y4yqmUMC8SlBV8d27w/fuBKER+lYS5uKK8u/uSr5BfIUukrMDpGkTVfQyHKih
fwYljMdS1mVtRG1oanh2dc816QU2Ex/d2oeXmHUsjkfyr0uQxLbbISlPf5vXD+lV
2DZpVKnW7i8QzEFz6Z8Q7XhjQfzD+qxGOhHhKUO8+t0VouzDYJhVsbET+7aM5iXE
WDnReGlwwQBqaOsDSuPxyNq9qt1eUYZl9eLM1AWey3h46Jh6fIoC9VdViqMNDpQ8
GbLTIm0WAqkooPWpuRWOehXC01U75zE6b6+ngDP2UNdqJE+byEu2UwGH4u2mtTo3
Oy0PCEKbAb+oalylWnHqXMzm7taGa+j1OoG5EFvz31mKhL5J6nD5bzV0vMWAy1lE
WtYdrjPr5aERaHFU4siTJix6HcaUKhlPWl13dQngbp9dJvYZyaKwj5ZFspcjwcNU
bP6GJdAg6nvPbasiB+k96QOgODN9yBDJlORgYJZ/ODqpFo1Zvxxsp0f5nvDZA5Rd
sjIMJekQahVAg26CeL7kdXvagtVaE9tB4Co02gaeqxi6wPlHG3c4tbUon/nS8KyQ
QRkxQhELvvAKdmwH5mSccFUazUk6KR4Wy6Tgygca1P9vkBKRUfVX8mN5e2v1vSn/
VmnSg/SfJHlgbH3pC0gKq+BIM0KwkveQHT7dvxb9TUOSXlGbaJ6qLI2z3dsK9Njh
3uoqnOJlnYg2IOK3ZQTy7vnNVpJ+iOvwSDnxUEIb5yXbrbKV2w4DMH0cyf9uEN40
hXXPNSgo9g3UBM0ogptzjZ8duuDOxXpnkBTy7N5F5FtdyZLSwIohfUQyW3oRinGm
8lo1hE/7uohLQqwes3l22SOMK0IaveZBWzW8jxu3PeSAbJKu9+/0qrDINP6rNV0F
5Dsrol7M+RQD80SZ9pxHwaS1NuejHGMLSb6gvXu8iyUBIrtD09LVfHxfK7bVccby
N6/QQSLbTH/g9VDmFI6Q9No7od4jysBosKE2yK06bjk7tOCyiG5azY3nvriKpMFV
syhjf/TD2qdpV1tUxG+yhGUyouk/+Hgk6pa04CKswlvwgYKnqg5+lPykOrgJNWAi
9dqLCwEmS72RVgqweExqtqMIXEVAYDJF9SIDc0J3J/dDgwEJO35Vc0CSNEOO+Luh
rxLvM5YDMgnN3VZuXWxUoYk9YsEGXOkqOrPw4djYyYyBOjWkURvyyB9VNBtu6aLj

//pragma protect end_data_block
//pragma protect digest_block
G0F/cZyRTp4dMjgN8FWx5s0ntKU=
//pragma protect end_digest_block
//pragma protect end_protected
