// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
matDEs84Iiju2moC9MjMB8ekc03bV4KVCkeTU4B5JLtabC1XLrIdN9+S1kqz3uqI3X7B+nFlUcZz
6HsF10aJFmUsa1ryvu5cPN5UrMDYUNSbVPiQCQZx8vvGPj8kberBd0laF1Loo9ZCsgtvK45Equj+
i5UjVbmJr4OC92mv/09onPoOL6u5whW599n8yi9C9o6BooJV6nkrrTU/dloEHToVhyovhTudQCi2
q0ZOddfzaRkV62dAkq5WJBAY+ZSnTL0vHB2CZzSu90kRCwEOzfnGVMU0/moKeiO6MZyhYNeEqzb3
WnQ6bJl+i+QtNTlpOx6KHyt28z6tVedwOyRGwQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
J89vmj1fcA1eKrtZ7I+/HqNc478XPlT42MRROW5XCidOvvJ0H2tdLWyV4efYfODUjLmYfH5zjgnl
7v3PCiyvB4a16ZepvIZhUkzoRAgkF81k6mAO6wWH23YjFuAMsumuM/jNXp9mVHdF54i2p4h7+hlt
IULZTs06fK28aE+/19ksOyd36ypZnj+GJROjjAVQDT6aBpSgOWSsCJb2QWH+TGOJMYflSIY2RCO0
0P8dqratA7wgpN3rQcaivLd2NqbVyeXW/aYUfHJR0DmBInBCd8I6Z7wUJHdkQ1YMXv1qb9rH5ikg
SunwwUybOixq2sa1eQunYLARTBiUNiuOoqKg+SUfa9YT9wU8U7shf7zR4IIP5cs4lGBY698dG31e
oSAv5at1kyoiLjySnS4UI54cEZC2bNNBMrH4gb2KAlDVJF++vbT0OAmWbSe8++es13usF6CHWkfX
o8qeFyq5ZTl96R50daJda43XPBsGbzWZ6HFleHumuTLv0p+5wArxZb6oQyQMJbYI2iIwXFoQXq77
l9UAvxr4DBpI/9GleqOGMNPSv2i4CvrpMOeYmg7fT4uMi6qGyIVMckrAw0bkUKDrc7gY9v2XDNQC
j5S+geGq0nLMn81S9t+fnVR4WQfmUFRZgy09XqIuqhscNJJzzOMIl1MyOBZ6e8QqyBTVLs3uso1u
TclQVckRERRuWfyoIhZiFqSB/mGhPdPKXx42wAuwJOWOcfttrsaXSoWGITGm1DJPVzMNY+LL1dOR
cOO51tcXGgFDXvswGPvxe/7ewNF5hZ+2udbKnMImAXG+veVFCYrfDl2Wt7ENkfD1UaIpdiEBcl86
zvJ0OOkq01EYUUD7PL9AFgR9txRoub5JhqbZZzgsZ7MmUMoFAdyqcVLwv5JJg/3qMRVVTwObjxAu
BzCVwZSZiuGlM3AYPlSGAClM/qC8xWAmwDpdzY1RKIIluNaO0DL5tLceU0SVJ+i3OAT2rDb0J7KH
/KsE3Md6GDvAD0Q75MDGRBU+CtQxWrippKp5y7I5Cr9oMW1WLcjQeqJZ6hZZ1hge7T2p+N7BgW0I
b+T91Gp9jkEEaidyo4PJUjI372shxc99pr4kLlrOEfHnjnkmQ3mLT2fedrtDwwvX79oo/LWP4r2w
0rV8CU7tDgIN7bN+PYA5D3r5WZdis6xElf2yVZG+1X3lopmLBBjeWV0R1EUpuhR6YGBd6DGiI558
GPXhntI+f6GxFW4L06uAPLaQQbW9fhPTXAVV9EBZ93u5hKr9wWxXwWqrRET3cSDpC6Z5mBCJEi/i
jqOprXQGQ8eiB7qHg3e4lsNEITuxJwEoJAcHXNebLBC+JAT0JAL/qwAMo3aTiydvOvwVKAQfkaOg
tF4GXZoptHeeqXvsGbUqbOx0n0x2VX/Tjrl1ZnyZ5czaGWGjnmK7mmgI7bN6TsErtGXXAzMlrFG6
iyJdi2q8EZGLKpAvCTcG1nQ+OcGZtVyTGoaqisHtuTCJ+ttsVq3LijH4p1wUS1BmgHhrAF/9PX44
Us/6jbpaBgJtnu12yVfXdCA0CF0EOp4QKEKEc2ri/+JwcwGP07ps5de+9WlbSkk8QvirzhF9BJ7Q
Eh0vtwN7H7Xtn0mSZPqSjXedssbh4qs5RQPT9qN2JaTLMvEK/7qMgF6oOXV8VijdH84JKvPuTG8d
9x7LVdJzAoXO6lxtRPziFGMTqzDxFqiocfyi/rXllYIVA3DwMBqwOPS4rQ5xEQXm67X7qbB5cXwK
CqR6arm3fsQqmqbXmpBsnZfwY6np8oGdFS+ZlksphMMP82vqAImWmzzX/ldktTEAyDovRhLPvANy
ABdMls+NzqbY/YXGdgHn1nzW5jAmC2cn7WdyKFJcxOzLAlFi8r2ALjlDMxIqQuSV63eoOxy2FL3q
FPJfNSAh9zN2jJBBxPaQVknrERSJXJF9ABP9KvfMW7B/kXJlV+ED1zI+UNaTiuCIugkNowv3rAak
NihoTbyFcomfZfpaWC/0MqCuLPKHb9mLF7VJQcLeGIx59MOHWluRIB9eKnE8RJ7e4Xt0uixPS+xC
qfme5UJXOVI8zBWQUxtk9GM0Jl0ta2Ll89YG+e9zr9ZVbcltSGqxTdF7VTkCuVtU60YxjRspe+a7
ABosxIdvASb2FfWAQG0C7/vR8a5+f4v2e11nmbV69KGPV+R7TVZbW0yNtJEF2gLjbHE/XO8ewBUJ
enyOEWhuQMuCkAphvGfrG/5xOpTfnBT/tjQ/tO/2lNw3KjXAdiqvyp9DaGqhPwPi+fKXdDaGR/2b
DyQtTgH3fneOZ8ensdp8U5OuScrQI1q75QBD6DjchxqNo1mTOSogql2S9kKOGgaEpoJkA9wzPlhK
uGglMMoRDqKDaWfrfH4ylq+osGte+QMwgv8ni7fgUoJeGdgDvYTTxhrEGje/ymA3WSXYcJmT3HWV
g/P2oi60oIjy+FuYYK5I8LcZ95wUaZCy0j5QtTC0d4XY+kGqCjNDIjPA9413xK10rpx3ZgCstQqy
GEx9A+4HrMLm5p3O7JL+QKeKG60kbeO19BPMJWyv/yGhYYIm+JK4JSM0Bn2qQz82Rweu9h03tZIk
WRsqMiHbKOrXgf7n90fcT52jYAUpgFCO/juWRJ79PEO08s7zPtlJ0cugll/0D4SuCRSVm7blixnE
gl/7ikxJVAWVZX0ZaVatb5OwcRDyBTPWwWRfZXpOL+h+O0NbBHGV5XjfzeYoMq3SaADdhGvpuRtb
jpzmOoLzQJEQm12TJm8vPX81U8zahyGPuD1NNxzkZzvNB8O8XqIC1TRYVw0227wonj8NIZ9PBm1P
v74vNzasBdohDB9WQnameVz97EGDe0cErG2vI1GdEyHjNUHKdZq8QWIUiFc/95YGH7vs9w7bELVx
sZeYA14ClDxu3Iaj5wi6sYm2wF4QhFjYCP709EoGS6cR4MVs4WZn1Zc0YgNd6MYzfYgF6VSFs4/F
axlzsY4h2GNaRLx7hPUOpFuCUrRVRfWi86+ujYy2jO8RQfzXmxqgcS5rcCyjeZ3DbzUzBZcf8PDv
pkVDJa9L25prO3UgmUHcTVZj/nfUmqGmoZ55GJfKOo6/Eg+uSMjcT9SiRiF6rz0KXYsuinyS2KCZ
y63zHM+RuLVJbnZhR/Uk6vMvvFc8CZbZt1gc6+3PWF3ymQ9hw48oCZmq3lgnPTe2rdUyXmXlbMjv
30zJZYVQBpGb1q5SzOgS6mraLe7ZJrCrqBFMfezOsufQF+yW/0dj/YTUtJSXUxPL3B4Gs2XtE5R+
17tNQYDY9509Gd0s7Mff0eIPSJ1KSOy0ck6VXgHfcgiwa5duCqZgwr0kioESnRjaiwoZG9hFhk0s
l0w+1JVJl9KuwuM1AqU8K79cEpF0Sc+2B9K84isQDv5JzmH4dtP3EYrFTnB7dZw2XudS60VbHQZm
FZ0OQjp56sXPyW/m1whn7tVnnai23yzBVYkjuQO9q5nlaCCyzCv8TllYOZ04mQcu0YNsxjBMQ3QP
3cNSwgPLNyFbzlNa9U4LthdccXYxLWB2I4kgRH5lMnTPHCqcxbjjQSP0yGoYHOGQzj1BQ6Jo/Tf3
v38L485mrE32E9ILrfZpEFNKpP4HEySpUU8qHDEIYqnMrRgt/+RsRNNuJKHmwWYffvoJnOyf2mzY
lINdhBgxRf9hJ7BwHLmg/dYao5TGkYT+kM49DuTIQmSgsNhEi02XwaaqMCfZ/zvQK+wVlQtXxmEs
MsW9CfP6Q9ruwC5FyA7pOa0BX860qwYzlzoLjROmfLOq3LEyWsmFPEtPWWY51eGnvqulNQvNU7Hd
6Jlv1bL8M+KnPnHTCE7C8OPW7MqOM7wgX4rLtxJOgJWNJ3lwYvxbZCxV0Q258rr/7luLXvOdOwcH
6gVS7fMmExu1VZkj46p/D0zWolxpAQ/V0kcoZmsplAUaEzEibMJW92l0xFMyQtpw2tVf6aYd2wbL
n4SmKgi8Ptqu4bRW0kMIDOrOjwiW6BhVWcCXHBU1CaiMUILXnt1hO7W1uZ+EVR24C8RZd7o6Bjzo
jSu5gp8qiBDf7NPxkxKtDW3icyffPtW6wX7DS2uKpjKDDA7P6shACHCPWAy9BNwoD1VAJ0tnMI0I
+0NcoITL+BuZF6tMARd3udup912MjKiSqS+xHUmvbqvOeRR2SGm9wW4V41Bqwrzl/yhRXHHZxFqc
26UfzX3wb1+ivpe9FgbAT4VvRtM7kT1ikSdYl5BePcX0gbxZhlNXCPvytiMq/FpTe/VZDeHMQIDM
x2UrQ/STsuamWEy4xEV9RNExbRHFt0lOXKngCw1P7EVPhOwIHTPv/00eaZcBd89OKRKx5XFCtJZg
kYAI/UHTdg1VlScEFVi0azQrD7yko849QM3rYMRE5vNRoklIlYHj282BJid7G4XaD1qW0dhaoriI
zGfWdImt0g7hRIsanN6ESa43m5VhFfZIIRsAEd9UvcWRVLbpyL6TuvdsIG8LefY2fA3oL91UYHip
zsPCcsKc1gWKj58fDdHGfFmkhyUjPwq9aEw2aFIAkX3t0iPJOKMyNh1Tok/l7MVpKKLlSJDmeJHL
zj7/scCRsonqlxHsHUXYYBVH5MLUSBkN2Uxc+RGod735tYsPoPrrv5wYejCoxm3YOXc0f/n9mMTs
SYKt8cGFaPQiNh+l4jWxl4IEolDKiFYEfrRulOYCyGePkmHZDgYXl3MNE+pwOjLTRMCYPPcjNKtI
2cOaog5IHAl6+nrAE6YWsKWWA3Jkil7C4Qk8xRO6tPQrQ4/i5IJhSh4yrjucowSVcQT6BnnneyhP
yMvRR2CrVq61IlxJ+V4qlny5bS4b6Ru6XOFw3uQ6gikWkjLkNdzITmGIAy2ewMD6eALf50NSDpz0
1DhGP92XLnj1tWuj+1k+Fn3RJr5t/wY6lj73VbUOrX3jY4D15V5yIUOup4RJvKYVuxiO9wsn3MkK
vUKkEQvA00jSVj9yQtxSLFPkSRpP/OIckPSenUPzgxVA/TRaayGJuZ0RU6LItasubDg4YmTaMb74
G/pNTCnlfCn60PtCcZilpI85iJ1KmMIWTSpY5qtE4j7/7HXeBOOlZLk9T8SaCZ71O1TOI3T6uSXR
DUoSjoYVKqzKA9J8htXVEobgupAhbDSU+dt5glpTR9TAwm1RhzTt3YpHER2sUl2B+radnwHv0qLr
t3KM+ii/ahKRdmwDuEz6FPJSrcCkoEAvDnS1VmdJpCu2/b+oUNB3rPhpbWpR+EWTNJnwgc/OTyya
ve9sUv8M1rKi+VoTqIJAfHGxhSvRbVgzk4Q4AWhIUyazSc/PaBXmHJl86lTR3tv6KeeDAB6yTB6G
JDNyEQQhC6EtrGYAIPA4TGLxO6KWb2OvPHq+6oW+WoBNQw8G4nw7Q0CVBVBTHmPFn00QYjBGbIT6
YdL4iuVk2KEYNIL0xtJ1mxZEf16rYBgqyvX0vHSZ7OnX+XF3axoO40VuFDC2MISfWiQNxZzdAckQ
4u1k/I75VS7WdWEq00eCfTYV6k5m8sK8me/Cnj8BJdhjELAF3cUftWz389c9NJq57NOaF/mmNJIm
Tu/sUQALMT/f3ZiUz0lE/BMTNVUEMS28T1aE6p8rtZfdBXIukjn/qddFdr/PZHrQOSF5/NVGuEri
DwdV/rEVZYoRJqR4LCe0QoidS5gP4kQdx2YGGiS0St3dfIfeVdVaGU0qHrXSeRRSPSPlSFy2KJKo
ABymvVmB0BmUGLAKTFnPnlyH3VF7y3JvQ2Tgm9cBZo9z6PDKmUNRsR0O7yMN6eq2bkQgj5J6MbAz
+K8whL/uqzkaupxmL9UMqXHN38AL8kfTRHniwnw9eMFI03O1cdjkv9LHAVTDBoXYSJ1uhYJUeD+L
97EeOLKyanfusH8Nf34IbFNgM+IZS60oqW6+K8eWl8/Hy8BYhY8otjDG2V2NIXadx/QDIPdfMUk6
r0QoXAgTodAxjP5cPoosJUNJvaNE39eTk8yFqiKty4KtrFv6629rKQseqtA4xGhI2DVGOQiuHosk
hNyF7EiRRyMyspykPhdN+bW4DcM56zo/80wRA5IFR34rGmL8RJgSsrqFBZRfH71tyw6+xY1wU+R0
JDHXtSY14C20885tqjbNQ65LtvmH8dcEXawD2uCmJ1mQaAW09/c36hqLQTJocpD02YQk7MMiW1L5
YPJX1D6rrMCWmKHwaxsVVtRuSmCREC0qyBykQHYH5QE9DrpVx4eQVZjun+Ytn+wKpCkeDs8qqH5c
aXI0/xzPz3MlfYEYfsUJj8h9kO3oP0OQR5jEc0Hnfhur/KzW8mDsFH/OxOcmEhQuYtZzo8PQI8FH
wZiK43aH2xNS+2NwXnXGPmCu+hMw1M1SDrwqz8xxrDFr9p9yXbdeKYxKVja7vvhSnNGnUi1OKG0j
P2uIby7txGH0ZC8rFgsBNEEh+UcxAaePIHEJxzHtxMcb84tBLW+jvH4L+M8DJOw87ouQmvoZcI/1
2y7QgJov3oCHq4TwlK0Ie1NwYiqMRntdgiJQfE/TBlssCoOjhK5yUYs9nIjo+t+DAU3JSWo7XA8Y
WfhJXuHNDCZZoNQOBLfxroCf84rucMSx9OS0N/4oG3EKJNqNU4SQSZtNRW7SAvvtYROv1/++WDTG
QFXTateHogzDCP1pN2M/G+allapDrwySaMmuy0tL8+DV51e46JVkMS8LDYcsb04IKLtdVtrwcFi2
OVGwFNv2g47GBkIydasD3tyUJfDeD8yfGbUGuo6qo95ptkCHmoR98DYEzspwiVB47KkN6LQxVYsH
Hmnay0OWaGzPRDHRX5MU7MXlyQU1W6XbPMX8yME6rMWJslQDQ667Px/TZ9tg+oyv0+l8O4pTLZNE
Pg0ISts8ikoHkh3cbxM0aFdpjg+dkkj82Ifm6QhAmMk1RftVpQ+Fc8Lgf7lV82Jxv5t7RqZBZCp+
Ls0lkwIxZ+glNd3U5Fk4XIS+jyV0RCMv2b9Goiyw4wUJWVpcsN+EHEdKZwQPpVGsBaB5Ibuc/bEe
A26Rea5UeCBPVWjeJanVCK06IE+5NDw2IyuJH5lPnPlt89LHbusOdBM3cWg2ydyjl7/VH2mTTRYu
hyAVrf0GwiAKaVdsGSvxrj8Xakkdi+AExWsszuXFnMR5o3cl/TCjJj412o/iebq/sLgWAMuvmYoX
I9ZuXpHrSFCpiEMZYTPZnWco2Tlrgvavsg8nhY/6monwlHx/qkMqQHKhmW053NdNnMMV+aVKTrGJ
wqvoLfUXMiw9Gl6KRpDQyRXwkHmlGB6AuyrUT88vpjWnUwPhExgYKCGweaQi4TofN0nTTe750Rpm
eHtZe33IGET91CbD39c+CGA/t63NVecWocpX/jVGa6s9wle6aF2xzCFSK70bBgbru8UPje5JhmAP
Yaj97LedJ6I3msCOozHswNq1g9k3n+BOElTw5+GbHtJLcgB+1j8hq5IrseEOa1pzgU4waeshfDm7
9p1TBi9wPmThNyQyCZ92iHv8gT3lFyglshmqrHp5Tzhfvmnv1R++Q+6/qzBvhfEgey8qe1apHLLH
sNHliTcu0KwDlfZ4rqPkiOLEy53FZeSDrtqbJ4N+Ul0H4jIEFrXmOEdqY0kOJqZzW8H2OmyhRFtT
z7SNoAL3CUjYe7G/Io//JWRiKXPORyIXOGuiwiwXkoGer95ynG5B+1c+IgLRQXJd1YkO+xpTTQP5
5mTR5ku3AZbrfG+PUgVHdjzJ+IvUjrTkWFyjDXItkLJHTSk2xMfDIS9HL2VkO4O00Fk13dLQrg1w
G4eBYyaJ1fRk3PasqhTsylNS9+DuWgBE7bTxJwOf4Ysy1+qDZS3/bFEUbph0jN6nTR8IQTiw4Dy8
NReWIX5VaZiDp/bSthfuf2wDjNZTHJAS9VlPsZWBpXmd+dYXM4gtkoEfRFI386NI/4ji1NklxZuB
j4PoOMvgSAhecl9+8ys5rD2OSdnXJsQGWHmFg00nk+ekqs6uglwsJHGMMsgLVNtXXH0cSHJUhts7
HIrqwchXUkZNDSQDnkh00N+nq1NSvhCXBBVRz8y1AGWeYiJe84VBFl9iGVd3vrEgPd0zMiWAFV4h
LrWqT6zYtwHkzBwUTvs4z1l/haxeC0yZp8vapAPNTZobUiOqgD5l5ZLMZlRYpECVcU62NILGSpmp
KBH5HHcA5K/UctISvN6QA1S2a0oYIWRX8iwcvnNkiA26MJ5ShrpMW/IZvqeNsU2rtR7rUmTp+cDe
N80Uoj8egGCYqpiVhd1CzzJ8c8MAo7LHuDTycnBv+vOVBxwENLjV4rABwW+eHxVF5Qh3b4Sz9c9p
fDRugcf2Utsv0hEPUPGiF7GjsrwXEt3IcPpgVjvBpkl+WsHyrdC8DRsG/btCtYaX2KobgpMcUwMf
soweLAXRNLuiBT58ymA7fVikl/2cd73/peuDphKyBtLfBPmWyJVtoevAc3ecyyHbS76MLLhdwj/B
7tXkqP9MZcuKkgXjPtHxc1F9PlAlhmjoxIuxfU8A1+KkzfwA1ArqhQgGeWxUJJ82SQhRB6wa6a+j
D7mJs/nafcxTU1oh1oOlYy3PQNSgLgqTKCbA+mwqpYytoUSaygDxsMxb26yfcw0A0Z4i3Vacxspb
+jEajG5n+Tgm2tMTPlExMkGOyH9xHG2LgYq2Cpgr9BQ7uM8I7H3th21xeLExufd8r46e+JbJuWmJ
RLBOlhG9KOeK4AFutVXcR4Ivx80RHfOMot7z1wFgskuJCqAN9WP+Coc7QhG7KruPfpSfgjLnw2Kw
1scNCHUWpj179USc6gxKwId9ETbwUe8BrCCMgYrXRid5ialqCvXuyJoAD+V4sJ/50fNuKFMyb4vH
lmh6jN3fDpYNQUFxPzLXnYGamt6YSBT0Sd+ndI7U2jWexw7q5gmtFzDssPw44/psuRb48UYWgt0H
LNMBdMtIh7DOQGKoo0ykbdUGpJmRdckvmxcaVipep6xejbrCou2jxYwBT7B563ONSnwpY41euU0p
X4O1mvOuC1QAJgzyqsRk4jQ3NLTQzVRPILs3+EYQrha0rG41Iv+NWGdtN/SECp6qPW24Vj0LRuu8
444Bwh1C38+Dl06XsNLRzk2bUFDz6GyhLamDkVAL+TR41TxAfhHuewO91p0ATlvRhDFbXtAn2Gwt
zWzGCD7ujEVM8hRHyxfrIQtaFesz2wM9RaOVtg0tBpgUxHeZy6LvmWvfPWcZlfsZMaiiLi4Ku29F
iobVjOVvGjlNSav57XPT7FA0IW3BNw4UBK0AkSs9B1nzNk2sFj8fzyU0Ldii6aZQ2/dNwd/Zlouq
ulOPQb4QAKoT+S/Og2gRLWXL7EKPbrtfyJtxbYHohOVJum0OyZpwvMK87gRn4nIHrJmNBzV6U81o
lgAzYsFX1iBSedBqYeLwRduIbuFXK+GDU8TErGLM+/zMiVz54ZpepwrKuETvK9bGLkjAaRZqDaGo
kb3gPP3P6wGUfLZkJ81H3QborgT93mbphEtvZzwTK+4OX6EyK1xKPaPZuoJAvuyyN2I2izbBJwu8
W9U9wIrjXJXJ36HG+JM+2NOmrmgQOafUeMlsVOPt90bcQmUWxSflhBj4MSxNNAVAut/6UmBRjUfY
Jn+m2kRQ02+8si076dcsr8MHPEq7gW/s39LUSMxF7W29+low2fUp61R8y0GIwqXbpBj3vNRPnH8N
kQKPh+7BtjaE3RGYkjuvUIqV6ytipj6s8Sfb2mbCVfgBKOkeWLkme3MBJJlDgb+jfaLdAbETR3cx
VAfO9atdDa0l7atwbXNubY/Zbt/fbSupdRaPdYSPWtgl0fgRL1daEuWmhU6FXNZAV2g+ZgEM7RNf
mapznTaBuc860+9K3lTMIS4Ho/FMTIFA9Fh2x0v8kpQL2M1jA/dC4yLYhslP5O06khrXFs38LqNx
jhwcYrqMGw8lDp94YrWF3ZGRyN8SrmGuxQgIuOfkncAsrRu5CyJpW4MN4XNtIqIYdnUT6c6ARtYh
iNpWVc/QiCAvIL36DeNVp9J2uLtoltaFBsyFN29cXWEloVjjsPpvJZ12Me83sdSSqACcwRK+jOg/
sI/R0m7iF4OJytpKzuv2jcPnG5NM2fmj9o3vhc64+DZmtwPAVU+t4gyKnWEbY3aVC2FfDkufhjDO
kuvaivF3RW8D/0WxOuCzWqtdxpez/yvWoxGybdHVGgL3u2eKAR5ONasPPkYru4kMXOlabcBQht3Z
hY7/1rIatCNjUWWLidN8aMBMhehG3LmOnoiuuufYPhmwI03PC+Z+eUJVzTOUAC5ozyYYE+h38PP3
+rQV538G+RlsVXU+yHO7iTt1ZT+ckaJvFT19kjAAshhpxF+cWn9rSkc8QUAvtygEC6vjaRabbIcY
+dgWHart4bseY8CdA2DzAEM79/U2e9oLqMPGo3w5hJTk9z5ef+3Mb3YMxOp3IH78SehFm4Jht+c7
nlOtCEvx7WD/49HZPIoDh3LSQ4JXCw/rrFLgXSVJ30DpbwDavM8WTzQRdAFioITnIIaZOf6nqizx
IwbuX59Wp3syo+rxzEWlck1LPcN0UsgUuxXNqvBehd+PkkaNRgldDGF9ekT1bhIQKZHiJM+8bto4
PdwDhAMX1M2uCpUDCyGmDs8kfCwgWqTmqKD9/tr+Zlg3XicQygyBl70g8jtse2gN7aUBRADNFMua
nOw/NWnwruWt99WH1HquW0Ct7UlInN2pj5UyuKgLhFfGjRQT6ZnVPnT8uSBtu+VyEmO4i3jg+h1O
ZqfGkDZtvRhu3dubkFV++KswlSaDYc0drFrI5Txyys+ilXGa/Gai/saX2H9nFk+hn5ckppebJixW
dzGjHVul1jLYssDnSSQyoP/3eKFHQOG2m4BtTczvCGKToIAF64yIwwCnse/hwvizFJJYMant6BkQ
4+ZYmFAnZuzHYARH8+5Gn3CCbTDaeJIDtUjkTBWc4rw1lj82Qe0xuCYQmu+uV+xINf0f5px4KqIc
GvZSRshavhK/QrEXuFQomUyUEaVp1DMLMOSHeNVCWBHF3UK6IfNSsleUmZLyClKDnvclaO+PVSOg
P8UmPYsvNoAt+Mk/b781easNR3vnoMTu9PsuOHGMJ3UiRJTyn3Q/wenQ4RIG0vRGmT0tzFViqskf
v8ile0Rux23O3K3kUu12uW2isz7zlfGSz3dOSygKVgnJ7BvevWZZ8oBr6CTMBwuhTV20PEZf6X92
V6YiQjQT+1aEXtzzElVLe7qoORQTYyTyqojVOGjtuEXO0AN8BMRe7qvVtUzRrjk5diTH6gs3p4WO
67MWLhn1Oo8OWzwVg30yIBjH7IFOARU/bmPuYcWv1GObLwF10UyqyjHA7PTjUDmgZDqgnIMQkpUe
yqOYQi6txfvqHhKhDFs2E3vUQ7DVdeB8O8ZEB+/BQRiXdtkQQqZ3wrjx19pfZ/6zUo34LlueS9hj
TmI36YjOimMPX1x36nF9ZMgVBWWWYX55fEOqE3KYNaItys44COp+UzThiS1iBgNBUAyN9Ap26hYm
U2bgVJz2kEDP6l0sILTNY1SGQBUSwu2Fmkuw3CTKelEZ3imyHxYHgyrYNU708C7UP00f/CqUmv/q
qjQuCOxs2Ds41d7hXByaRRi7uX4adsRgkQ0ywq5qXci765hJ8mieomsPF6M65hTv5zVkIhxwrLtP
SwrkF90ebf1zTg7LHVOnT1QuV87xKoalCbMAjZ158L+JIuVAE1jw0zQrRfCwx5BYwvPmXKGg4sEb
k0flfRG5cZytRH6UV9Zs1SrV4GaDCcinDdCOgA57enCDy0UndBTkwW6ZHPOJJDRmU0m19Bx695Xb
fK0JIGYtKoMkFQWw/rzYT8YjrkNY45z9NitARMs0jhjNBuRZyCFxGqzXJd7pOBT3CZ9jHnN3EAg8
E9+E3xnUwB0MuIBKglhWJwr71BWgBCqu+P+Hp+EzoQUbwI4GTLdzF8MiXAfjIeoRP+Du/x8YgZjl
BVGlnU/+Jc8nLpsfI0DaoU93ERYQR5VeCcwJglVidIWmmYjgQfbq3Wt4tzJr5X7SH33vRgFeyYtL
GMpDZdXXUn2vwfg3LqLS9wVmlMgS5zcacXcnoSQa2Dz9EZUvkowCytcPMxsyfHiPTAaYFvz8YA3J
PIN5ABemoB/YabUl+0gQ1vxXPvoGQFE4bn8AXcyqKvx0vqeXBgCZopMQdAHHLqdf3hVW0FqduOc5
A/Qu23SQPCGNulZLsuJBQlmiQzpTpqtBuHuCoWiFj+keNLi47MdQJ0Bw8j2H8QXiOKhQLRDZTFfb
DZWNQ1VOmEzYL0+CY2GVtNLTgPxMpcQdPhfS+O7mKLm6h7mL9iblNeqkTe7eW1ipDXTNBeu+nQGB
9Km3ROO5sGpN7tMcX/ETgWZBipq4hMdODKxVz9Pq432YzLl3muh5Xop8ZO6oeiL1NJ+BglzN3nRY
O/ISUKaJrOGWeGd6S0rnPjYWGaTzdV8mgJgI1RZZzZp8q+T+GnNu41Qoud+xLyiMkI8UbZkPh+UC
jFhcYOzfkewSpgs40OIpt52hImOAg8mLkjARw3SSkN/vi06UdbbgvgbSKGE4FnGNvFTaUmKrMxYl
S7u3sWbxPACHBbHVHODfr+emd7oNBqa7ixS7+TdhjnnE4GM3GbjYfDK/I0w9d63w9pJu9+DTfhyJ
x16ctYzmt6RoIrTcn+D2U1DhLVFp4jHmm8tSCovsch8x7jveuMlNzSK4P2VzkqYxBGNxkf28u9Kf
q1cNu5Pfqc2GEy3M+n5nsq+vAbiIqVV/M3Tn4rRf+cc9d4kps0OQ757Bth44Zet0mlKfUmx/y+la
EtxMPcS44V5fLmBM829QBbV/ttOcFZhA8HfQ0bJkcPreT0/P0xOFX+HpxVzhO8PCOUUehu2tRE/Z
pCgc7+TlwwvzS//8mxHAOsTtetF52s769KRtEYEcCCpLFNurg7/gY9Iq4L+VhnusXfYrN/hivhwp
5Q2/lYQbeDwse/V9bYD9P/vXKENFJSdP8bFHyLo2TDMQtHNAvLuusRqbUK/B5KPfoJyh4/o1DNVs
Sr52R6c4gcRi3y/5haXS1T0dpnAIPpDJOsHvc9MVCNdBIwlm7I1EddQ8QHk8QPig/OzC1pEulPG0
g/VzYRJBB8uH6kSkUkkGjkqrzeCE0PfaLolYjazcBol+5IWVfJSIhPka/OjJA3zkIPjaxlbsTlap
A3n+3RfkT47yDKvkR7zeNnzVhQSGl0Cc9aPj3iSVMg9wIQlsaEa/6NiwConMqzXf/53G4mAK8Vf4
1msxgoCA6bIC22svIGb85gQ2StVtJNeotsOsVjk1g9+95eJtaurK7BeZ1OZo09MejAwUTHryIKzB
0IgSETLotPM69tf+SrtB7sJmoFHDcbeT88n/uXwyuN+2oKcFGdstaQL/OcaoC1gGBB0eL4zLp0lY
2jSEELHQSFD1KhBnPAQ8VUjweYlywOm8HkCQAmDyF5MMz1geIM/8gSEtWrRkNKKc8mcqCSlpIsw8
SzU5s0pDTBscLZy6aHK4VPPj3on67rZx6Wy0AAIoEhi13A5Er4A/eLRksrUJif2NaQHwcmdf5Io9
aBM+rcBWT9Al8l3fOarb8HymbPLbI6OCN4LkLuLRAisfnMMtWjd0NiLRdl+FC2y4+nmAdgWu2sTA
3ScgRHPODD24HEveRXMpH6KmcEkOdS/KjAfLE2EPUuQTu0opZz1Ym/ENk6SmuUp8oDWmZ2RAlGW6
jXgWhdAB2eOGgbXaWTYMM8paJjPOl2hSUp8AEsg4K9AZ0cEXb+uznHRTc6V7GFfxQrYxo3Cewc/G
bW2B0o2+eJzbw56Y2m/s6Swwhd720n8Qjf43KwqPb7z/KyGAUWq31Virz94GN6O4jIFfUAotPpna
7gi0zNhPkgynMMnreA3WV0YzpUY3vkrwH+FEtYPmkdgGMsI7Fq05xEb0IEKht+hGe1qIRFY0KoEk
GWnSzBsAjzYA9YajazjesYvaaXLGoZoxvxfOhASxWzCzcAm/ZhCKXWsgBz2WxWep4MtwAXej9/H4
rJ4l0KICYpjWbfypSpcoxc9vCV3myuoLC4jWuxcW1Y7xiCC9XsDH5DrBw5zZVe1FQ+YzRGbe/GI6
sMA948L40ALH8hqtsr7ScCAfhaX4ZaFV4tcAg2vk4a8Ab+Z3nQ24gB22hVkZbvh1KsODqo0wxJKT
qVgEo9MCFIejwphktXCEY5lH2kUJlg0JZuukwMP8y/NuaxUUtNpJ4Sqwy2o0NPUNxFEvkce3xw8R
iKdkvwKYYHqnR4k+BGSCb9e2BBIButZB5ag2a4QjHitQ90GhaFiCfqXNw1Ja+Sh/fh+PDSNey5co
IFmiMBN7KZexqRhzDP51S7/nyjocCKEXBLMG07lZK9ehTusLftkMiF/rBrytXwc1gF3DFu4qM3HT
u4oCc1kMDd0T68gskQKza8aQ5Q+rC/bwAuFEa+MobKbsmvEMdDCHJX/pOkJoOCfg9g25W9pNYXJa
4uqBbtWvMlcVJDszsCsr0rKFjIF5GvC+atCdkpxoGoTjQ2a/Rs8CYuBvqal1ivWM8cTpp6mFCD8e
AXgmkzd6VfrZgM8LS2UMIStr3Pijael++dXxhokEAHfKrJMPSl3CFwfZwP8S5EurVmWVnwlM28vk
jk8nvjOsSsKdapXPwu16oMntt8cavQzc48IxI6RgBCDWstMeMA9JI2GEbap9EB0PvOM5AO8vMM64
+bC7N0gNvcy5nABhmIpIvS/TnDBfLT5rU8PbvsCffvcv31Y1kHCEuCDicR51xiA3UjOQrN/aFYbe
YH7RF4VHJN8N2ufv5PkkDgUvOMN39Ba2WdKlzJCPPWpFNh0N7/OaykFN8u5L5zjrR1+QOmbuRDOf
ZPdtrWskdGkbAOH2UU8dVSnwmfQgJq0l3Zhaz8To6HWfoxGXBf8HoP8c/ZefSazefqhn8BbBK9ru
12mHwLYf14tzdszZd7VfE89HF/DDQTZQym9X08+A8bowmFlIBRED6oglunbfry18BF0qzN/0a2bs
mYzHcQNpNmpCOAYbtuHmuIAERFB4DTuvv/BhJPCzjpPN8rRfELk1NUYOXTVMFjXgg2R+uQOqYonx
wu4AkXBTr16X002reHh/JFOhSat8mtDUxTkOw/ZLoqS1JUIjT1pvUDqMWV6AdkM3HZPaNhXQkxoX
JFxHyI7mmgh37m/NpGYQyt319H99ealedDSLfvdqEZS7A09kWof8M6/NROIf5ju087tNtcAWzfGQ
5owAKi5pj5ZGSWno9D29V/xeuvv85V9WEEaf6BKbtprnyvnSdqxzPl0kR1sfOJ3NfVrkwHs+gJWG
/Y2pM7w0csEL71GlE4XQCRrV8glaHBBjCcBw8f2wrfEiwKlQmGEydPeP9AbWehfCqBuAkWF9y+u2
yOoOlSXne+OTleYPMqUxObHbFwhWxd5suoFKU2WbjAKjN8gYSO8y+hzg2Zrl3rM/bOik4MJiSPPJ
nca/1yL87Lcnqp8F+No63MK9/Kd2rc0FHTCcA7v+7/3JgDIOSfxFfJ3B44P2mdOi41XhPpnAc3nH
KgDONSzJcdiw9Ffaqi8McBgCMnMB7LGr3PJfF3B1UAK2Pq2RLT2aCTuyueVQL9Wr8nNDWWFj1e2X
nXBOrvMbJmkSiWUMbghJlIsQ2RISmdtN1meGaEhGg7aK0jSATG2dfPqZ7nec7urVp8Lm2tKNN4M+
SHA76Eh/CZ3Mnr3I+H9z+F4BX5moR8o0CxkLGjd+IUGCjPZRhagRZC/r5LqMbcXfQIOOOpT60iQK
wPi+Xdftmb8XkAXKN3J3YyMSE3/YEDHmiBjie3RkHpWlbapmuw/BX/LlyKW+84oE74tdJ510pvS9
fi8SLEgfP9da/1A1UvykASiFAO/VIHbHyeRVpXbakklfY+dA1lHlCftCKV5k7WbWuwQ/izkFhqr0
5Ca9hhY1VJkcYhhIRJdPf7qdrkHyDUO37aZ48lyuffbbD4jtLVM/+cXHJRobCYfb3ndpL9xSgjWr
otbaOZAbnqot2OtuoNpo+UsZAiuBbvNwmcGoA4IR18VStBDf/3/Gzznd3Gufxk0D/tuypVcsSlQn
7BcMZf6kt3Ji3mTKb5NCo7yBTPhu83l3pyVbF0mUCMyDMnm3s3bQDwixLdpWL+1tuhJKJpXm21Dd
wX63c4k+HyD4cTXstD0UQdphv07hmeMI2IvQp//dG3dRk7w1Pz+Uf8dSABE9Wj8vtWPtvpxg5qZJ
ZdMthgV4VNOYYnFMxfabbxT8TaS9DDSdOcmfUIBRRIeUhoNXZz/H5UDfyLvvV3ayLCnCnjiGGBFo
BqSUFVLcH02lXsgLtUcAvJdr2MrfLlfoNvVjLArg5mLp9C6fsOs9OxqxdzzxasdlecfQmzI2nwN7
Yv4/E5KfGZtpSvTaZRJ78np0DcihatWoEeroXGP8GE481lraaq+z9KtRHOVWl53J8nHbcjO7q7yn
ZdS1x0Cl0brsTMiCGAJro3eoLL28kHXNX0MoESNn8WuYtzA4d4CBf/UIiPzdW9eZHDg81IkJDi6f
Zyxte5jeg8IRleyNZQrX8mFbt2DLj+tyFJJzvsprWWjYmJGqMyUsVx1dzOjmv18I25WIhuvYdodp
zpPZY2aAVztgjgZjIKgA0EsTLezZBtRUcpTryTs5d0JU48nU0W26Kev2FCK54TfGGVhCpXGboNTr
B7QLx6yiY+t4pdc8Pxu0kCXeP2848HvLM0Vfj5jlGuBUFMtGeRGcMHRThkZDiy19lQxENE6Uao/4
+Z2aHlCBNDaLvmv8Y5SOfCx/HFR/Oly0LHPdLgkQToaTtOwKiVHZj5NxlsGZY5SXxSP3WwJRivoP
WwbHb6dlyL0PsCipW7oV5k8FlR2gCR3hQ0i24KmlmtXea93dOpBx+yYVDmwyUyRiaijlYGPMnUdy
Q40JIpgq7wMyMeB9mq/+ULx7sqowa5XfiazmsBg4OcWvGVzd3s4fj+gSQz9CK6PUcWTkW7mdpGlN
pPJVk1PzmJ3uWpcO7N/Tx1wIHaiPsYDIl1He4/cl7UbrpQqXN23Xd4HuIO/UzG9JWEC6OX4cIaE4
TcA27PyKXmnm4BPbNyjqA42+cf6QXKuIZLTlv7354aiNvUH4+ipPbKFnuSdfcKf2YDetnlQwR+vG
vhWSLs2uTWAFjQuVY4lKQnN/YmiHLA/RSz9wHULT2iP7VbfaZt4nTDEThvz+4IU8LrMT/DbHFIAK
IEclLsfDHhZJJp++WuMh/HS9VQnKplVBCkYg3nFgtOdm+o4/skHtuXJk9n7AXYKP7C+f3//EyhDO
s8bkL++06oIk/vlu28UtmkigbA3o334n/7th0v3A7zgcTbepWEUH2u05sV4fu/+OA4t4L2HW9/Uz
8KVpk5iUkO+LC6YKEXlwBuDXtf8aIqTy5ahf2rX0ztYndRH9MMnPl3bNMs7deoHzdFWypgY3uV7M
a+3bgtylTWeY1h+eRHsyEbQk6WqMi5c6CdvWS9c6TrmkjEnxQFuz8FezegzZV5ra7cup3nbUQKsv
4cwUJi8s794mfvKwJ/oJQ9wXibIS7eJD4xvYgNnxUHEbllMsohEE2sbF7xHRc2ugLxbpBLDkyhsd
ihTdw+RlhOPndkZnBL3bX//1Omqzc1opghxznHgw+qwo07tozng/SWDLrDCtKyAc9ru1yPexsw9T
Fh/vL1jP/e0u5RUtuOie6xNCCHo5+bjDB3AJURWw2WXLc6QXDTcil0PjAn5hEryTrXNacQwQ/knF
FckDdKoqS1rRXShtlu7n1WGmUUSeHBrylxAcL7qWx/YHgbFS3aR90WlS6O0GkW11ZEawMJNp5R+p
8RPTMW2MDBDxxvO+UdFoqj2KUkiCP6HsHtIt1yRA3Ji5gRPkqvEGxTUJBo5WuPEAxmVA1Nz6ZjkM
oK33e97LEPdi/YYR9lTs7vRwMj4LrE/FyUXaDjbJn/tICITGsRhwS0o4J4DRoXK1TfBuWCjjG+/A
+/+cWga72peD3x0dOGnurIpyaKDJ4kiWlm0t3pPJXwa8OyFtAd7Qo2/s17QyyoqBEJ7yC59TI8Eu
pLSgDF8QaA9o6t+Q35uZ3YH2jXjWOpZPfMjYb0D2yE2Rsp0s7qBuExQyuMfpNS6TY0ViuDfnJmcX
NFXvshXEx2NJjPOtQW1FQYLT7twE0f6Q2p01ESM9LR3zAlGLn2ACSSVqAdwnfuURgAaG3tHOQ1fn
EVsiyIxJDh44TJHhMzKJbxrXOduZRFY/BNoWcPr8qEBR9/Xi5xmp0oL+iq0T5IiJ8tQwW1arn1Rh
HiLOL2t9uSGb2EIGTy5NfPmvte+bDK5lSnqTvb9c4e+BlliQj6oPK3PqlwGghK1RburVB2AkTcri
dtN3NE5pt2JynaUNaeMVepO44uePYiH7B+Kr95NJ4mxzjOED6takglfLy85odIil2i5nuIV5vrm1
9qDJljtWuUePB9FSMXuSr8ktrCTh2NABVhje1F0xG9P3a4gAojAhNjx7e2VdWMyTjGvYTLXBH70J
mRkeB6+42ugjbtRlpvjWlkmLXpFRCQzg7qCWJ0yurMDvNPGuW95QHTYUWoaAUI9n1AvnlutobO9H
eMbLNiC3DzqDD/qnQyv1HeEzhtEWRE1STfPOSMWtKHm5/xIV6RI9HvcAph2fSM5hieJNFV3XzXNU
zkywORF/wbNxumi3Y8EbC2tpHR2ohLZGlaVkTB9y5ZYgfJeXxQ4gdrzyaOfv2vj5x54E5/BH4owS
SH9IRpytHxQptXw+qlhv9Nbnd8/oSTKDPOHsZc8bJwKRu3EEW+DfeRum0tlZHbKG0weEY9n/dA8R
dTzmJGTHa1Y6y11xwAmmd8RWMa01Vb6+GPaJlZJ7bpyv3S0Rqi4UeP7JbhvcqYk/FEk99h7qoJlY
x62uUwwFFtcUo7aSyrpvHfZWghiKiG5H8Fifa2OK/d0mh+y8vlebuR3y0AR2ngdix+Y+jITz7lv/
AFqTHacxNT00bVP2wa6oQJvd/Jh+Bndx6kkcFH1YuAbPnvzGcXPI/ydzVY+rBk7xLdmuvfaeL79I
8kOZcSfV4Gw+N6OiBdsDh3K9fo9+uXYid3WqFszlBMCJ1go4rc+0YJd+tgJAxqZmYN2fjB2vOep/
jpQGmIIdArbrLOxthNIt3+UHkFI+3wrIgcv0Pc51vuA8cgM/behTuz7KV/fntIQFPa4ih9P/0rEC
BFSwkpwnLxMNWuiZVovNAx2jLNEAFjdLbeW1WrSIUh0d8ZnxbmXzk+88AqzBvRjhJRl+ZVePuJJW
uXA4btCoK375vftyfCAbiOiXzKNiwREOu+jfGscR+NX2ejXrERnWjbZ1FDUW6zGiYVMnaPU9FP8P
aQXncYZJgoZGeiofsAx12Mu1zERu6Tw2vyY4MKAJnwLvvn3gB+BR+j38GprUfjxXdtWbPHQ8PaEQ
m+amcgnwBW7v+NLjgSZqmvmFT/Rvp8NhJZMC85Ii9MTj0A3HFL7p6mQCbKQPWbhwQZVocdIowcXX
3ANDxR0mgrVN45CcNHM0WWej9oI4KRwx22BD8vxyhetsD3KvXt9Dlj0BwgLRtsw7jpZKdQoAyHkb
zRH9yRmmF7elfvyYcsukuKuFHZkgcyX6YYDe2Ah4A0UGctmj83hzRg0EHi7WOI5NpvRG7FphGt4b
87nUauM3Re+hHLwqbSXo9eK2l5Pkq9XlPAJqXZpe2pfJs/7P4ca1cNQn4vlgYE3UDl8PcYL5AY8Z
thv+TSmsUSseaP29kOy/oJk/skliBMkvmdBZGAeWa2CskSXknAJXufeoEzru7LuOinjIiMO7849B
cjAFTnXh0uPUqUv3ULcHsjYyVLTQt0KqpgW6pSSEbwYXbdHux9weokHrpsRbwv1/qgzBPNi1A5Gz
tF0F2pjatIFRVME2pFsHLQG+XNdn1uQBEbl962kR7THAJAxgE6TQXsdnD7u1YU1b8YB/OmtKAemn
YMtx85/VXxGPKuRfhlNMUnJ6puFuK0NgAmFu+2dHcnIVB2HJnajVfVvx5nHujoithcl2lDP4eC11
tLTj26mdowgH9tQ+H8wO2enUUG7DBn44eFgGQlrZzjVLAMndxILbwHRPYOlfva9LObL4E++Y0kt9
2f7QB7MIKY78HiIeYt90RtpFKwJkpn0SjanTim3ptaNtv55FOk8Ko58QX7ChPNxyYO++2yZpXhUX
ZCIAts3kipDnUVNdgJ3fHnIi3137pO4hzVwJgVJplRu1BpM2RIXgFfkEF/g96gs2ulWKOCbBX2Q2
TtAzWBJC5kwyINSJ6qs9MoTRSmOtC4U0G/kf1lejV4JrexhbLokx+TzGiSio3QGB+fdaIcsbBVFD
2VNg1A+0Wvgqm5ZJ7d/1JrZp9uRmmU2526yYWNUGNPO4rpmiVom9LOlgRweqTxEgYWfmrYbLEvkE
ZjS0tUg55peBKmJ435oBPRpf+4iNq6L1+UJlxRf88/ARwxA3pZw0QrvBHVBjdgH2gRpg6T1n45Ia
GpheAZe3c+pQQUajoCBJRKJ+kBMrBvDbk9zFNYfkXhtxXKiq3A8XEgSZP95DXSPXh1IysCyaIJyp
moe4z+pBB93Lwty3Gns7eIkbw+PWy7Wf4SxIJNc/RnAo4w9zVCmrPnKAGU/ZkP+hZVwQ837pHBkW
9s401qbw/F26K74hyVZCYNlTi+ASogBGdK3dIhPuhogUKfZa7iNAp1MvPUYy/lkGhWdft3gjqsaj
Ec0LEeAQezl62QzmCjs8r7uVLskq3LyzpPSjHb4fPbzKX/xMTt2ITxhu4OysDyawJDbvWq+kM5dK
cHZTx4cxD/kgNLQjweZel8TlGX0W2PrUoSGgESnsRR/hhUHwCBGoXwCJjlymvDF8lX1gVtsshddb
TQr0x/7ZK34OPXbZD31oQhgs3rcyi8SWl3vON/o+Qkv1pDPEDgoEaz7x7Qw+q5YwY69LRjIMc2Ax
Ps/33X43v4iKHMlnFqN/Ay+GTPTD44QrfZlfXsX9zzSNDHgSMi1RdxKFSyMDVOKeMs1mYHf1G+M2
Neqa4pZNyDpEKYinDT8UxnRP8uwCr5TzT6FsnrqVFBJA6FnEhupaOm+f4KwhlzoZhZ0G1ADmDr47
8WjDGOOIN22gz4ytj2cJA2YiYwRKYHs3eHeXfvMd5/CNg+7groHRxIs5ngT6ZaDd3RAHt9MBTGi1
MmobrH+RPBhE7PsKAZSmqJGxdjcr4HFUSCbYqgZ/3yQSU0HEvekAXWwhveniRKBjwKVYFIzWjAiL
AVjTjriBiH32vCYa5ZWICedI8OqQ08lP3c+IOtsqcoTUGmBZXWXffPejWXdSbBFWf0YGo0Ru1z0f
0hHgVNBmxF6Sp8v88P+jo0vECQtHtAoLkTK4WaGYSZD75IjQU3EEQr33ymz8DudkNcBFPPXBgpE4
SGhxxEcNAvY57h8QIyjpWxlFwwl3AiU7ltiLJJP3MIcgLjOwsj302zIz9iYFqYXqemQzpeKn3jga
YwS2L2s55SYLyKAZprbqcN2FAttkQ+1DWEdY3Mv3/KbNrZbeNbVMbGMX1ZenEXs7Luu6LtkriImG
dzkroW2N0hyBE0QKijs7A8Qa0ZROW9kfNwt+/8LnkR78QEPWYxCyJbi81w8Y4sbkmW5dwqLN8h8A
x9IcbJV20yzGL5b5KNTUvieWFVamy+oowKRzKM7PE9O9AdYDTPl/5lhxjaDDIn7EFy3qrgFQpIZI
jvUQN/sXZ2wuubByblnRHEZWVu+mDfrPPsXukctZU+HL38b/xebd4b5yRACFzJB0fV8inio2j/xI
ADbyY5NYb4yy/DgDw49kEvODXP6t/jWuHL2wMjQQvhy0+WvtYFsmGWJpTkPjRpS8sUCLVkI3l86n
yNlaTv+YZWFca1P9i47H+Qsy1eo6VHL9Mdb3qT05Hs8L08d7TwgczjtsdA/iOz4iy34+LvGfBV78
6NxUcHsKm5tUpJttAN5tcU3ppF21n/+cOwP9FJOVGVb3mWYzyUJF1mDCYdsw7IEuWQswMp2i72V/
csxs9ZyxuHEJblWGVZ8Vzajfyfc0xFu6yeJQtDq7BPXhA2m4g2oBgKtRqvxlDptOn2H5PwIFa1yI
rl8B+QOing58fKjRGMvYZZlclVQYdtcNQVRV6X/8ER9xTtTj/hSlzjkcPWapmjw8bqIYUy5KwSX+
wAg1kaySsJgtcwfOj+YnAMHprWopDYVVqtv4R4LoQ9H2a0bjhDmRZksZ15MtM8RgfZJmAGOa9Oc5
kwh9B4l5bEwVVhw3s835cSUYf42U29msfL3kCTjvGjzeq/Cui5LYi9NcDm9UesBCCTIX0U6XQpq+
4IiaYfWDrAFLk1NJI0rbx/jQW7YxVD6EFGjAYXvYcthmH9LDSyoJTcfV/Gp0Ugpo0V5I4NYZPJJx
uchmHrDNSaUyjbq3zEF7yM25gGkGSb+wIyKXb9jxKjKVpRIrYM22Os91fzdtzD4vnj8jh7+j8IO7
3SbyIXCRJuf23JxshYP8sfrXJl9xePVPUV6HZ40Zo0SrDraZeWEBI6vS9iKzJ5hu3fAXwNVGSCxT
1r3zczAneeK2csx3zgGpDEIBvaqVHrtGqwh+3IxNoMYxqBdoMYGxTiQ5oSjYFz5lj77nYtV1vsT8
ZX3Uzu2JzvDCu5+QOybZ6ZDdZWPIXoN9HFK0+EfykOqP6/FPPBRxTEOntqciVCWVUzXGKZr2ZLb+
BDEs9KvuItnQX4OnpFgOyWQ2XkP2LvR+mtfM9SywEm2PVhci8q1NhuMsb1fKnH+2WhA0WNFqquHX
27E1NEFFICdfA/Uj/q/1/8xAR8GbCY/6joTv+p4mdEH8YJjampTLCLPSBq4V7U6IMDRAJPztkf/7
2SmOyCk8bnuhH+/vQ8SW+Y5Wnf0hrh3AtvhsaL7ICgTgQDFrBPxdkw7dl0ld/P3l/BtpZXqDnvfv
fgmG4qaCIXz0WJcZkonRWm0DEOcYDtDbqS9lJnpQaETIsP9NwnPAECgFE9xNt3pAirN15zvtWclL
fgOhJaDN/lmDoRSkJMFwcv0J4Sj+Y12ekEhIgQdMNV5ZZq67mQefVbV+to3DNfiHobLF8c31S9vt
CS9V/n2yiq340wPC0QZyJ+rrqCpfPVaHkn6Ujwc3fQDt9p3MdGaJkV/nNwjcvDuj/lYq9wyEgGc3
ipohGx3+/fDL2i6Uyapt9BnJOAlr1sshhntXcmkDh1bQ+/bxFZGjbj5WvXZ6nL+vc1f/uCVQ2umD
y3BMTTANzApUqOQHmkmJTRDYCBdEssfidnrVo5/1tr5TJVMZIl7Tz6w9jmAm9CSgAC7SkYqE+QyA
5Zk4GitAA8EB5jG1MME0L8FPg0A6YDO/+MnuoUY8Qilcgbrcgwd/dliFmucZTje0b4ZHHr5iECWN
/iwXnGJ0UWNwsW6UaLpVwurn20oAtrkMj3camJVuIHK2vlR0214DpyDl4Py8Z4BAcp2YOb5Jx2N+
2C7JUpRCv93BxiuAWCxL4bamB97OA97W3d98QQc5GI1Ic8ZFvCqemWPkvcr9Bdka/xmajtmiIPyX
b0HdNzwABn9WQnr3vTrMNARG54fzFelf74HX3ikq1Qem5VnXotVfxpw62t1R4c2TR4sxlCUbA1Gh
6B5QUJswZkQLusxiKhMpEkIemHhhJYwbVC7MUy2WpYOtu8dS6d3l+0BDKKuZj4dDjaNKqFx45yE7
yNJx55M5pyVlvj/ALGgWcI6UCvqZXVZSszsaR+Ffm388CdR1K0d1+JRdBDMO/NNgDIcLtdOxdKZv
KkQMoSiFNMV5N8NcIKUlSGBF6Z0P5UWzRLL/WeVg9gqtQNS3cx8kMd7dAj/mR8yU4g3MU6n5fIT/
cV6jQ6otenE0eG6zWfQUcji+Usn5/kzzERCl+NM6+bqTcC3wa2NRU1THGXehKyLShB9pgXrE1KR6
e3844kFgh73xLqjZ5B8y6xN0t6u1w1+i3jQeERIMbIxzZEP5SxaSuCBoAaadyqjtT5dX/FLwxBKs
z8/shzTZeB8MryOhWviOFguqJr/ZY/mDEpO18UBVaChiBTAbm0BaTmjzmGAzqltHHukkga5qGm1d
XkO3SrN7ehdzJTkHROFSTQ28kdsIqavWM27C1+aS3hSMY5L1ms8EZuCwYMPrR51XR/fDmQIwblqD
Sfuun1bCbSBIRDtGHiRJAS8Qwp4B2ZGyzubq/UdfA+9l1Wzv1ah3d0Qda+y/CT3h0EftTiTGMF+s
xeUGIpsJXxtwlwg9gWy2OAXa0cBx0Ttur23YtZL7E1ap1NLDgpj0KZxJGCifr1l5oqEXMRDGhKvd
EhkxFJ8/6hG84s+5Nun920y+c/AWgRwHrs3pKOUJYHXY5u+TXIssZBDhUSnNV8Q9+7rkioxEGxx7
/ns3EGBD0uqw35RopIkHbhDD+PjW/DOgWl6WQSfXSlXxPDCY3BY3Rrke4EDLrQf4lPaGhu61LeDn
ovqLu8hBkTauRK+rY9rVLy5LwlPeUbah6iJJuaTNrphvbCT/MRPcoFsV0mkDm9jApOuZU9ahyjQK
zo78/O6rDMoxx1FYxP65EdPUsMGDzOlHKMaFmJsnYV6I36QfWMvJLKFNG9K2fDuP++qAdIBwgK2y
NxIyfPBlBCGywDs7JZUbA+SGUF44l2zv+A00EnI9LHcFqBMpJYli/Yh/9N7zc5AZj2iuqie4f6WH
RVNZAQiKORkCrf9Y4DDHEg+9hqZr4KqbJCJEUjBt7k6WTG61v5+UvdEqZw/76Zr5YFfyHx3wMWhA
uByjO73JXA9godUJ0xM/ZWuH6vH+gZkYbeQs5gfm24ffKLFjpvyWX/NNEvBla1Rl+EvNka2ydftS
ZY6j1ij2LkJvJ5qjxFr2lgAWLVZ/fL2I9xlxk48Bx6oWeYk72ixHpWmrBiNAMvQ0YBGz2zp1ak+I
5W55NwA4jzMBlYExi3UO7cn8+f47itcI9Klrx4YHLrKPgSqVXNGUX8oVzKdVzCweOk3hNP56/hBA
OO+/UKGTcNQY8n3UoOEQ9fNGwOhYe47ivvcpLAU1xUw1vh8zwHaikyvF4/NafNTKn1KQ7bReKO4J
Az4/IwDGFg3FanBz2jxFZMAqRnOyiASCYMoOHuNK+jTnfPsM1KPWXARMDBaMvHjXpz3qzt3weN5A
TtjT+DgiTh3LQgTTMo3rt2AXkv9oHpgX80xIwjeaH84A7mAAwb6zr64CFP+Bl5SYEwP5w8kK38cV
7a+GfSvPpY/SLwcnWOPc34YQB7skJk/PJhxTl2gU9uTExNhaW8uQ6ITdPbTK+KBmBJLJzJlSkUrn
QEy9U+Inbm9gCa4TmtDAjZ7fyrch8N7wF2N3TNtr7B3XHyVeYvqFY1Q8xDnmfYQWJwB1SBE8Zbgq
NyiBrtmat987iunbtTthjn63Qw6293LEWi2MQnHSZUOyLthOOIzzinasznfpOb9lnjgF9E7X3xfJ
m9dEyLb0nBHJkXog0AtxI3ZH584nlk6AeoUr37WYX5pj/Deehp07GkDb+a4fgOOXcOC2frtrkvCc
DIgyQSIORWBswjJHLpwSdEy6PCb/f9y6ZhOj0HM3ZfyecSftlUdqGd1RaQR1JBXJX/4W4iLzbVYw
r5Rk/Thzt344nW1+1qILm2J3INFDC2q3tkVuhVMZcTR9sxyscXb3VDhCbziJTwhj7prdl2P/6LM4
LOoenzYiVK0oLvXPtAA0Ysyq6BhGrcw7p798xc7+koBauyJJfjCxZe1bwRou0e3BbhQqNxsxRiOy
trEj0KYurCnHKJ1bECMfW4QZYCRF2W7drwh500jezn+vx6WmLFKSmrZJ7TfhY9h4IgHK+gVWq6rw
5aU2zs0bl+Ya1KK6W4JavhAe0ycbX1cJh7NRSl7G3JwFcPLdQf04MLYSHnA4MfU1xqeEMl8s+F54
+gwvnOxxy8ae8ilOTzyZqbRbxk0NAw65r7goZZrTNFclrCgHeYjWe/54H9BkgeS2jl4DbRjSnABt
35796pLNqp07liuIBUVCGSaH49DY1PfriGaiR+q9xLBTMi1ad3lVvZFLwk6KrYndLEiEIhbTqGlh
ATMbFUIROPleZz9/mdcJKySDEAqVHfBk0MwbUVpnYq/NZLvv29amANBhLH1pfQpikQdxadVPoe35
GJQ1A+0khoiGHPyeqMg4FLW1dyTpvGC2hOy9i41zxL+yM24w+co9qfZPIMJ3iQf5HVtYMUjxrcBA
X640m+nUKgzdTFlwXw4QOjobdzT4J97cpbtmYkbEjRsm5xg8HoMpG26aWPM0PbgPt2ho0EmX/4cE
KQuCOB183BYnRAJcQGjA0eSchvGm5OzzRbT+7w/Jq4xTZGmI3ed+4sDXlUPqVMOxmkJ+41iQXS1p
9PiH8+yMkw6fa0Mnkn6D0dxSEV67WEMsPmtsDhyN1Fs4Gn/BmFNxEy21U8GUnJ1gbs+1neCzjCTK
PjHab2Hcs/AdKHdI4tn8Jht/2w9elb7xpv5ENfkIrsEPYEM5VNZcNed0UZpVluk2Uu87L9hnDln0
QC9RaFwkGqN/FwRY8XKCfveNxlQjEFY/ZncwX3O5GkUfyiifjhbbhnX/dDS8Ig5fiqvVRGsLPwbr
lCJ8rr+w+iT8GpH1zprWb3ZJga+0TwycQpPnx/jtQ04Tbv1WD7wJa7FKkvH6VA7IVfezp2oGeape
rYeQ3GzlN1XNjydjhy1YSfgBI4mF0j0Sv9EBABF81bRwHD4vmLDny4L7JWMq45YuND5Woa9rlTjx
DBPmiz7O4qo6Kyd9l5jLuzritUhmvnjzrAYns5o9ldeLHig+g3dkozP3eSSLtcCNPPqJZJp3C2Ij
oDHE5ejz5x6lAS6ztBWdyd7feIXLJd5/h8e02MTLeaT/CYim+CUOL1alZw0xPNa3+0YUQcdoTxGW
pCU/y4YQL8MUSHmEm7Xn+g0pbiKxXHa7FYhhwsqVpeSaRco5btarcWtZwiPU7vEwBnCt++aSY3Zu
VdmxWPk1HPHh0BxKkOduhF9J0iPf146eT1Dw/n72DevES3AmxPfPSuXFjeEq2yEa/tlV+2o5rDeV
1MGLRfZ7/ECizQwJ5sX2lXupWGe8MLvWXPrWDyZcfCHVcdOGGb9fKp4SJmUZdVC+JAHAygikn9sl
9H/Rxv1iOrt8JsiC6h52+Df0PUDt7vDmAF+WySbzI+SOh1pPTWx2TaM6jgEdrPBs3uTUQttJFj6G
XLUQbZ4OGYPV2pw9XV7+zy3ElnyNb6luLIcRQFStsjFm54j/TOe0ussWem4G6sIgMbpc17+TZ9Kj
NXCB1mV8HK25K0HTiovHV6mhmTa7ueJpBUGYhw6rJvI2W2FsngOu+dBEVufF2yUII7XyMd0p0kJP
FR2WUMupqmO4miA/cM30DJ9bu701GrLK5KmqqpSinGGwhDoW2XQDZ4guIvRitiEQKO/fQkO8/tZG
KkbZI2t7w+0q3AtugKZ0DW5RglkTBcheefiBI+joY0DJqHKzm0XOptVu9YKn971P55rKTY7RzkY2
KtIErHvBzUUEKsibSKJkt+8RQuiDwVll7V1GANAnzKO8O4ORLGAfCsduQSSk14dSvNqs7dHZJI9K
cXGhpxZ605EhegZEwgV+rnr0r+6fzHtPopezTcIri5f+uXa/DM6w+Itr0pxn5WFYOkR4J59Pzrlh
tmpcqcE9j/zgTkjmHA8FvKQhnuMd8Nne7mFGpNqCzdcxxMJ2nlnPMdCgi+dJFYprp4GLMYcRuGL4
fqLniiCizgpP7Un5bG0xmZnhbVDPWg4o7pj5uisZQJIUUivVSmEhOT5RIWmFkqIp5bPvqbAi9gNT
GpJ/8LZxXJ/PiFu7cFVdyRRkRj7/PC05h/141Z5lWTf4sSZfP7V0d7xhPuBIOXWaLM65W9W7GPpx
Ogt2STmjcdagq/dXsE8yrOtodGq6BvbqB3ZOnibaA4l/PsRTAEk29eInwIZBjfOQppXnwL+dvbON
1FO6oTg77l/lVTqP3m6NHcN4OIl3fPK8hb3G/cbam+uQYG0olPUjRQVyg6PVMh3JGoDu8kU2Twxj
njSdAeW3ZmIt3z1zOYkF6QoaDY1V10iOXzdMNQKtHhUx4vUze8Xuw6IR0MNToyFLb4KBQzV5SfKW
NMkVlGaLGmBJX3Lze6C9D0DjkRPc3hMc+UjMmNDlrDar9bqIBX5ce1l1MN6r+LwvRNC+V/EuP9qJ
rjEpVkOwR4+joIKrCPDmggctj/vAx0rq8S0dck0CmVFjmwqV03QgyzBQl6u1OdgS5HfA7DhDK8+/
TXUsEYAWiFy+hJl9LSbBi8vDaxmmL0x1AzG8ODdKIjf8dS9/feR34hV3b5ekjEWav8ElnKdQt7Sq
36zlj7xzMAGeI8mfvgtSzwKOcZEIi1BI1DK+Q9h2MFlv4qgPfeI+gWYIkxzx9YkyQijrMcGeKsYO
Btj40Q2ehfYSUjsvxUo7b8NZV1BIi3xqKjJ9h3w6mBbiate/Mpq9AnCf6sIG4t3Opmtnpyd6cQmh
YhiHS2J2XBoqoECMHTGezd8Grx+7p20tafw/ZiZoRrShVXdLBjVG+7pX8Iob2jCsWQ73CAS4GK2t
G3S7Tv3oQ1QXy10FU+B44hXX0inAc67OTW5l22yxxR03nZ0mctf/uJgTz+sfSlGL5UZZgxSWBzUS
SFB4z/gS+PGJwGP9oy8EjK3VrTTpKMJVo2Se66QXO/Oy9w6ckwZpBNqvLQfc7S4+M8zk7je+fvic
2/qUKzAVSgVGT/mAPbGVoTuW/4ZIscrmv0JAtbcS0RVtPd8MFeaXeSn9zlOeaBfTvbZ3giLk9CjG
Km89D4T1Zsl9ajQB8mBYJcDrB/vIyGdoUhWCSARkz1y3UxrvBMGnsQXCzjQEZOSLK5mVFpHHdhGb
NQo73O5ugrunIWDnPLzVRSCr6UBMGAG8KUChvw4T7qlLoEctQQYj3cHobqF7CW9kyEN2vNewsT69
+yqZ6MEz+yEoVNp9CYGhvGIXjpC7Ldw+uNNEwioKoAiDBtRnnLvajuXg5zHc1v23hPeGsvZa/TWf
oXFu2FKXvrO6n11bj94UejTp9BrdPwsQt9b/JDh9HZ2WGz/W5ZP/cfQrzLrY86wybXCj1izHD5jR
1N+bDulVDFRyuokGdeXHFeNMKKiMm3ge1YCm5ZbyStCeH40PZsiV67+Ej8pyR++LsQUDhwuzVXFd
AKBWFRafMKR8qJhifF0TPqimNto7Fw1Ags7zhaDkrzrcX3oeaxnyuHCzN2YdrybOMXrT1TW978pE
RGt1H+7iixBeyycQCMjqnYssdtfLbbvfbvZSwsjuM7HZySXJ9G8NktSY1XXx/GxIn3ZScfePsSaA
YRLArSW+jn8haE4qpBtmr+S3+3G8bGuAvMcdMbcF6t1R8sX8wRqOTn35HEEumC4IpQ/0KqlzVM3r
MQGn4dbOtV9N0in3oo6LQ6/SRotuprDKMdnK8Sri/77OTbL+8xfrhK4K0eUZ3U5mMvsaA4se8zS/
aI/TRaJGXD0o3xw3eaYxJcf/VwFWWQYHdKE5eCEP7qlUwAgd0dhr8ell4W1XIOE+tumCt9eR1cfm
TB+2H1UYFyCUSv4yUoQ9TAOE5agU/mCc1+oPjGaLHs+qzR6gIw8w/ueWGdrUwSfz0Ex8J6crJwOv
1u0vbUOfRxksGolple5m8jlfDgakjoZV9T7tiRQZZPnl0uscF1jkoCDAw0aOu80mVIw0/+hGhUmh
KoTxCngwi3I5V+kSAwthB9HMxXAcU6+dl90Pw6h6NyxR6NhlNngOUKiqi+83EJT5YRRNY186Lvx6
ilfTEjkjn6vkcga3R1wAHXqm+2s6MBC15RckkaRU+E40vPM5fP6NAA6m5R9awSgMguJAUJ26VhSX
kfKGBdmFSAbr2la+RaSN9PEeqJU9J0e2IFz/fBHz5m02oyuGoDBuLp3vLvJTZT5psKzGcbfjS4W/
Zp+Y0Yeb7TIzK9nOAXknsTLl73jFie6tpdLqfoEUw+0FYogtoPnAJaIerSk8i1sQB1GxaIQzpaoA
IIVW0MaZMdRlwm6sdjbbAuGC+uD92iT/tuvtwP29jHLY3+Zq0/W5xEK/Uwqzn89Ma9hNKqk4hpeq
tIvRo+XELQMABhBRAHDJGveRRfrW0GqoRQz0RV2vlOO2t12EqWSGYkOWtEeEHEAsRoSqkg7Ofl4s
vBDi2AC0xYa0yodi1K8TnBojUaBzXF/c5kn4ljjujNowpfAV4KwCYmO2LnfGkBHJ7sa9llOskP6V
rJYEIrAQZsi8+pxfFYRgnyzNJB6I0RDYTOqWXOb6J2KDlTdUXznzjgo8JMPE0EWbDLzrdKe0GkbZ
9Zlq2I4udXZ/iewaKbcgGLI7ajNuIIuJgKnxkOVK7dlfURc30is5ZsgPq3H37vMWO/kze0egmO4Z
NFSzj27KT73i7qnFNQDFlqIOB1scCEzCER84NRHteiFN4IrAwyR2YH4XT3jN4DwQwzFeE6LOSkec
GWWXGilSQomS9OOQKMBJ2WN8x2I62YFl1J7e6P9b9MJTaGA8kiLUXz2ZoEmQGYSefLXQggpIgx8y
2E9W7wlcuR6vXN+sMGHhQfwL8/ibhrimksk4ukySb5P4lEgf+88au1+s//18jvdVY5VWleaOXuhF
ABo+DejjDq3A0UwAZvJow+zaJR2hL5aOXVOQJD6g4q2j1x506ObBQnQygZx1+rDd5unVrxjplU/Z
DR6GSjQQapyWmYSlwG6hSst3u2UDf9f7i5S5FiyjxucDvoF2Z8RSus7H57d3Te1RmQ43mQH25BO+
lnBmgshrzpfgRnNrUr9GDpYmkXeqfgdZaxxLxTokK1TRlAQXkS3zyROyvJz9YNlx3bG1WAWjZUZw
H1iq/AbKw4/XdT5AcuHk/iJAnBMKwzks3WFT2/yzjr6V2Uulxcw3YwaJiSATur7i9GHJCpTGlDfN
zR2i0b8AotgRWwtW2snQx9wPhnSFgpFgpfOYTXJu8+d1oCoQyehqF9rJgC5YOGIjXMqKHLNHdYcx
kLqdN3hg72FsC9MEPnvydQAYcPWuW0PAw6BeHAiORfPNJ8NT0A2MMRYoMLsDviEq7++yph1SGVRn
VTFapDLARA8PlJ2jQZMTqAQUyLITJCEKNzsHbd0UovvOa+Tgz+OHOmSW4S5jICQJNlPNR8aCz3t/
r0FgWDKAy0RzuffwLdAumVUd9DptrAxBo9OVxkp/KfJzy/dZWywOI5Lp7oR6k/zLCZyMn6/NlZCu
qxXjOLtPFrQsCuI7fXA/b/mY5IcCg5SbuE3NYAnb2ok3sPyi4PWGXoUXzzB5c4DrvVOOez4XMJuj
ZDyePbdUdAIfcRlXAaZd2kh4OHh+GoLjfkDmo4uCrscbHwOMGc7lkRzF7AJyKyhSQwcfMpAl6nqP
0V3HIyNMXtdrdOrH1XJbMREcITBiO4jxiX0VBIo3d6IwVfwmri00p3U5EwQ6rLXrz1M9zbJZPVMt
mXxVV0zZ9wrzyLLkz9J+W15WuRloBVB8/q7/qSvzrkm+oC3y+8pVfeVG+8OXnTol1BmZbuhMA2oT
s1JaXoZG/2M4nbWVm074+HLf3ZBNoXdoimSJqarxXpjo9MjqCvC1VFjWlO30VZ/2a4PhidkC+arU
zrH4G04uOU3HjcLj4dedqKfBAO8zTprL/WUKTWZEh03VXhWOpaPGM2DS7SqhKVXFd9L2SN10K7Kz
sQKGMmmmeDFTC2KqZEKlAccNtpqrjQcXhug/aTONv1jVDAfIw83HpAThaRnBvYosao0vqEsdPVCA
sHULyaPHmDvFgAamMHs3SPx9M+8umOaC0kVFWI0t9VDFvPlpcCnbY3h3uHTBumphnNN5CpOnjISO
843ypAz6BvcV0WgyMG6WZMLpJfTq2wKhhL6XDUBX3CP2V8LQ8QBmstsG7KwFGP6v1ZzftJHWAJ4I
4SigpRJF8teSMJemRhGXQeo6BWsC0ZxECozk5jJ5PJKXRWbnDY0rrzR2arSXf2ho0bS3SXIDU2oh
wdRdE20vXaC2yJe9FULPzIrHG1/gC1AY6wMQ28B8IAk4oHnu7OLIquMAjFYzhnZG3VmbwHDxAmjF
qqDcG7mX92AeIuA9fN9jw4VRMRvd2YhcVOgEEr+PdPfPaQGWKkTO2NURRe9XQNvgQ330Hzovs2l4
ZVfw+5AQVt0mUPEm/WaYETmHmbrzUl/rbmOiqMpxFvHQAmjHtOGYSef20Z1MhRpANTUjuz5kShEY
HmWe0WNWTmFyVAv7Dn7RYUzl3EypUWdg8SusVU9jF5D+++BacvxSyI+7Ppykqpj2W7TpgWnkqUSY
E9jqCuD5F2lofLanRhwq5UOIgei6/E36PACn35U4EMkjFCmDOq5/oncNwGlem5sxK3+uv7J17zdP
1VtetgG6EIrg0udJSCZIAswxEQdOE32PeK6UaV5L/QT2hmi6GWWOSonUl2Mn3eTMaP9qRVQKb/Wc
3Crj2ZnfEiPWqWLJksriPTxy/08sS3HZXPUAPRnuZ1WYtyq044Itd1MgeFT019+0RPjjujFNahmY
Xl3JzmQQR7YSF3SuFqus7RZcww27CzpALH+Gwmeg85zu1afT28rqNgOA1DHF9GEwTkKmBKps80ZV
RrzJP7McvTbwu7FYpMdTqJG+w9PlcagufQfsKPY0zXUd/Oe5dW9L7zivaOjI+ma/ZI9AwO/DplOO
HmBITVg1p+1WPO+eAxGXqX/LkwBbJSfZzBGn6OpASrVRhVwlt+cqqsEsVpNBdFfXrF/iAwUmnviU
Z4f9zTPRNK/WuyUYuqjYaNo7wlIkM8ks17EzMC/GuQo/B2m13wzpyi3OrOS+w30IHVXzWnHg/Pro
kXqt9D/buBWp9AvJ6J/r/SuomMqEfIPjd8VxHXiwFmyyzlmsZKe1cy3ZzOYJ+iStHhwfQLdW+3lY
u5IrjE+VUjMNXdm16oWcl7p+Cha6eCVd0zy2mOmUmVryDsj/qQdA8IVuHwPxnTfgqiwbOm4Z7WSw
UT7FyKUhcIBu8pF6kHttcWlYeoCoAv+CvC1uioT1JU/2I3JfyvHyMTFVn2ZoklQ78XrT+UKKPfN7
MchxyQ/l+uxClRST66cmsALFQutW+dmSCEIixhEoDE1NU4NdyVD0oGQa/H0HB62U+1J/m6FpyvTn
LZQq5UKlW8yQbQh0MTztKmpxAHPRCdkj7JavbCq4VK1S2v3XC/8ef1K/aqGAgLZgmla4aGb2CPFN
M8Hm9huI7xdULgEXGn//Lk86x8Ssj64nRCeFH4ZMk7ZG7uUIj5CQnu30oNIp9w75Q9vxUzcLls8D
Xfun4f8wvBnteCNIaf5okm9wkfjiUnces09AhxYwI9DbZ1MlgDL0OGMc4ffoUFfPY9Sxl+qXog0d
9NR+7oZrOLawUVHQ9iR2qr+PzoErcrRS0ZYmbpE2AglgMQb2VHYmmBrII7rpzQJ6BBWL+PUv7qfX
P6Z9r/gQQfrZiqZQHgBRPErMoiDuAwXZPRtTxiRGsshpyuMJ4LrfPeB4+BI891xHqLdKP6ng0+3n
xLbS1HqF63wfDZ/NjSKMrhz52BsTS6XOjvCqI+20TLWaPw3/mbgmxrP7DX7btTqCRtHJP3erE68F
93iq9cnFPpMePCdOeK0tSrgyQTfR82rXI8ZQbgDpKAzcHYg6kicupRL2CC9MJD0AR9tFE1t+L+uA
Qu9Ri7r4/C1ICCGMu6tVSgK0O2B2FXbrjT0EpChvEg1iM3G9onwJYvBmt6sxxwCFA24Tttw6e2zD
UF7kbmKBGk5NlCFTquSoHQfzg1mIyT0yrrte+KQGtcTxYxRx7/qJ0tWw762onUeLTBVnUqQXgx41
jzwNFBg6qz/hkkPgG1A7b+cSeHX7MQpCXCx0PWeGL2qugDq9G5Fp/pS/192chBhbtPEt9gNxspWW
o/I0BUfK7R6D8Yra7xN0acmloQokef7iziicBUaJjzvLEPmZ891yqtycFhR+mekZa3+ZWxeBgTNz
OSsRm5SONtt26TRBw+rEOEfMfKPUE5y7HeotT0hZ/mSjVx2w7XNdK0QpNKC8Sw16ULXmNQgLZENW
yKSkDTVJwN4BwM3ozMIJu1XLMFu/gMLvTlRvtAuvuS7brhgV0CNxFioeYf3fyuNULi6H22qLTbs3
UsNWjfnry1SXlYJpTlEn26ILydLbpUzpu1nESUoW/o9omFMXLQL+atyNOh3XX/2rytIN5xYt4rcd
c+yhHNURXlKsg69aN/MD7Ra/M0WiiPZ0/2VZxPRI99KpjbYrn6R/nAwkUGh7bI8CPsF8Uo2g3R0o
SPeK6gvwz/rqMjxNynlQixEuuxdBvU5PG1Y/zdTILWez0zDnrLOGYzJeKMdiiYm+GsS4pb7YYCC0
ZWzPwzvpYIUfpdXiBTl23iwX0NnKyQALHahhlE92ILWhCMAN7e6ObTuFcMARN4X4rNxLxuZ4EG4S
OcXwOIfDWFQYhIW0ZZ16eBnHoBgfbGrik3kaDyHf4SaUtNXglxJEvA10qIjY4zdc8fPPo8LU65ys
0B+nPjzvSrpr4djDxpiQ3KPrcSmZE8ue+efaSYv9wtHu3+z0LRTAv9juHCmdZberLQ96azajOL46
Bd3qmaRlfHsyi15Ry0UQD04nwANP/UqPNSron7ni9Gow1oE9HxIbQ/HXiVqM7CHLlMBpKEJZSbjp
Mv6h1fp0IhhhxoXq1bxLqweopW9s8PiGFlU3q6iMDvC2701iRo1m3RM7SEwcmGZE8T/1bGfPr4Wx
81Q3U26t17SA+KPFZwvpQopdxVwm6Nk2IOJFdRGkUYxpBZnGHYTUDjEbRY4S4hjJ5TzrSsatnkI1
PkDt82sTp39jWd5OnlF6ibIDdO4mfbg2UdhpkXTX8spEcbzkYN9XnqBbXJjOfeap+uuZ7zetjUhq
u6BUiZ3dnKXfJ2wPa8zUiDb3Z89S7XYNG5j5MJqbxLLxLN5QoAJwOgNn22v2Dbrio6uhPRhSJf9T
wzN3cm7x9cnqSwFeRmZqW4bNuVsrYOCULUkyphqFOb3LxlATaAzn8hidwPY3trJY05wsHeo9KZoo
nDsRDmklRaoz5UPjFZ2oKot1EzKqJoujx+nxZgR6lYRpcsDNZmDV/htFZPmEKP7zT8HhUZ646DXb
VZvTK1zu0d2Jaw7OxkWwe/7YivviWxB/TikoVR1clv8rwcw3z+pPWeaUpr1RdvLAo506lvORe68W
ckxyaBetnkbXeC56wTN8tu6P9ZCm1+FfdwIttJksyvXavdJqnEoACruAW8maFK+Zj3pt2dOFiX4R
2R6beMadkXCWnZ0HoSO52Jt2Q9hPebxsAJ3loU8QA2BHz2EtN1Z/VEJL0GRbWR4GYlDEsGuvSqT7
c+Mna7AmTLDpSJyB/DONYzZwVbQDF4K5kUmK/mfqHEkSyfywSiUXeOspR2Vq1B2V7IVpp0yHDJmL
7V0eRe/MAzsYYjNAD29p+kr0giqkAv4vqaZza2Ckikau3fByFbnedImzX7mJGhtOKNjZ727OMrA9
O03W8o8a/FnMfujyDVtByVPSOV8ZpyGa9gsG9HztnOZ00DIZwFnb6XUc1UTwhmDWikjF9qs5d3SS
gwRkX8wmgstWyJ/V13+cXZCeU6SwPsi/XpSJzx2mzfqXAdksF2mAfOQUCuRgmibdi1CO28jIacyu
5h3UOMLwfXjuc2mM7yk1W7kXVkskmx18izXbYflz4HtFIoYUecfiEteoMMRiA2EnMtFyEsm2Iba4
EHwI0BblPgLMCHpgMo89iCuNGtWx3mHTT2EhrQ9hxqMNiN11Xf5Z35xro4QfG1k4APpYJZ1Fvmnc
sZ1LRzVxuRc0RJov8m2+oaMlPSr1rK0xB4p7h6V2/wbdFgMa6oQgjm9MOTd/9Azottu3jrcQxnqB
5JES584I8/+64Zxsi/WLFRGCSUn3ZZM0KRgwX6nxGWiHgkf1gGKvmabaUUUyBTgf6t33IyVYfSvw
bI7ZsNME1h7EYvF6q1VMCNTUgmyfHuoblb0IgeGv6qPDJWTdjd6PmcO1p3+RWJCvDG6yGwAzOlzi
WfBzf3FfJfgFrsWKNArV04T/BDlBWnLJ4KJZl7vKdtpp1X7GYx9CjCBE346pWgCUuwnUUhix7bfC
X8OG0G8QdXp49NXm6XKdCsL0ADn91gdrMwutyI0lAzl5tC/gKxpLAGYNApBgNutW9RH6SJcndTB7
wgSggOFDpmMZ+OGqyNX8HwzMd+XaBG+hNpPop4P9q9XKKpz1l/OrWr9unEE8TgmsISsGSKfQ6rIr
jRUWiwSdbRFECqcxWROHOJbPxDRBVQP8BgWo4pVt0PH1VyTJXXVvuCuMakG0AvttSSRbYEUqKTGv
MT9t/PrURJm+nAMj67YGlDT5y8h2tdjBolY2iCA8pJnzvu37F0N716zo0CAX6aTSldSHoQmKWSp2
nqhcpxiT1upxbo2aC7qploaVtU+JqVG3e8y6ydqOmPIw5zU0pgiY8TVYPuhXvjy7OzVY9VkLxFUz
kTOkSXruRhTLBjbT7VPrCyIZ3TeAkYaadbyDKd7khr5Fh+lhFcemidCsJJBGypkEt7Yh5NM4llVJ
6o0O3s79hbcAgNd2wFa1S+nKFQxj0q5cHy7y4CL6AsVBfNxmTwv/ITB9n7tea+GS/zCjRjAlaUWg
TSnlxJ64/5A/ve/cezlzDsapSxmalUX76hG+j7cuFO6AMyT6SzMUka6t+TTQ16jv+R/VMCqfDnru
5ag+gorN6PNzQ32GEJxBPm2UR9Ozpi9Z3/j9PYz8P/KQrPXV8LMoYz3fC4ZgHyZsR1qQA+tiPxar
iy6tbHfQNzQxk47pqNpoIhs7Hl5f6v0Y1Ow8fBtVHFgsfHa/PqWJrl9nMn9wqHMX+koLUyMMKjlq
rK68nH/hIhtzDJ/ZRqjJ/imiJgOf9RF84XShhz+e7nOIkDf746GwWqn30G1xoQC34ffEUxhz1F7e
ttzyiRShWLamoZqloQlFPRhpWUDMFprfE3BX+YYIhqZMGdcVCPSVwllwDG6q764WtS1RRdzC0+Ah
FqUMOZHBur6UiIetR3HnZN0Kno6s+Vi06aL/E06wB2umg3eovlCJkvtRBPn9SrOmscQ4FoDoZ+NA
LA==
`pragma protect end_protected
