// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
GnbC9/lUW4FXMKIMEItDL29ta/8VxtADYRk2ucvukU5hlwE03rkmHA5MmJmVnHgT
cvliusGIn67oMlgdEIVGXA+p+qgQ2bg9MqgyDRiTOwVdfQM0nPDjV74f75Z2yp1g
ykPc5GXY4L91JJP+44GeRN6j1qv+DEXNQjjPnP8t978sQkPNrBA4Ug==
//pragma protect end_key_block
//pragma protect digest_block
bq103nyGFgpEenEkqSAbVP2JVcg=
//pragma protect end_digest_block
//pragma protect data_block
6tPP1qyiRSZGVjl0Z3yKSkMORuWs29xZuRGPaHjryKiv4Mj2goovHUVi1TCEtFBo
WDwO6A9n1l66mRsxLcRlTK5zJMyA1zm5PHw3RnJTEyYAy5RV9DTIuqnghoAifckR
4E3+WVGbODPBmySjQ/LPePdf1tz3IUKTMBtXOkhztwyANgVK/alfu+g2Py3pKkUu
7b9Ax5n/y/wJaiNxbCG09OlpIgPTjKKPNFddzomf9krfyWmd2nVAli9VEbCVeMK+
eW5V8BM35YqukfPAWuRxMjnPqbmQ9/30h3LCysEXgSDlALqr/ZgLBj/hafLdGjvG
26Rk2RNiq5vnhRT7ZEV+Zw/I1NM7hCbxR+sIjvMsiGPzKxImbvqnSHw5jhVYUNKR
2qUBz48K3C5XJ+St9PE3IIs3GW2sETIEKp30uhOeujHYrUfYTmo69w/dPG38lU72
RVugyZK0lVWxfNU/zfKcyYIHseR8WQN0eumWKEFzFYnJYVHCYhcToivuXPzun6/q
m441R/QjiCnXGCP3fvJOoI6VdWnXkbrUgSfmxpnk5xKKsWbX1p4u3tl31unsW+9+
vh6Nd8jSmupFsPVEuvxSehlAajQE1rsQEUJXT58Y9/qbz+k+eG10nsmM1fCjPRIE
upBlGRrzGuluKpq7kiNlX0fHpUjkNdsC3XvIzVPqxlx18aAfvAJ46A0/EQdG53j/
0HZXVGtcMTIQz0/z4BgfmMwvo8GkN1Bp7MrSb67RHDwx3Z6DAqaNMOVtps4D4dw8
7GwojVcWk4MykE1lKSZhNrZs9jCvZxGP+6dxq1t/Xrjo2iECozpG3IE76Vuaqw5M
XLK1mudJHQyvTGmlNri++/6Zsi/cGBxr54c2K7tBZJhdcAXLzApliQHPsMJYDG96
t8SdBwqRoIEz8Hny9tky8DXKST032PKx7drUzSNnwyMP13nPLt3RGL2MoioPO6rx
fGK5qklPOrxHBvB5jjqhh3BAeeIDiplluuaB6ft9Fs8wLTVbUmQG+21McAvZdW/P
jmAv2zFhDTzXWYGpTXSUzJ0jbaf1uKrx5AIkeLUsYml5QnJvRVa9px9BAEN4JZIr
SeceR8u+icr+KRqraDObk2FSXb7xSe+mR/ZqrLjZHzSXfiwEqWT7X1gWZdRG6bSb
B1teOdbjbJsb4f3YIPUaN0P9TyGAiDy857zZUdvIjTN5QuiTyt7spvmV6x1qKvcP
MplTkZX2TOlHAuWDwrIk9GpNjXjnMrMVxbQkLveQ4ns+Lh1EPfVLvw3djpvGq3Xg
D3ASSexAyygIYtmMDGiam1ZcpLD4RguEi54P6bOnP9apV/0bwB1trmEj+VrpER3j
FyAJ+8pX4oaP2dyAfaTZZUdEmw17x6sjNuBQa7ZLJ7cG38dYMIWntB7UUoI4HT4S
llTgxda+qdnyHDx9ubiEhybKfms85VXWQOeeq56ZidlYKi4890m+F5I+A+WVQEi2
bann/Grkg6xdBEkVb7zWMG7PnVoGwAFvr2hkYOf+Pq3S2KOpTYjaq4O9ej7OwDS6
BSl1iv/1jnippY9QvEW4ESTfJiDjYgb245ltmvqtrREtqL5QFNnMWlPJrShgEWKJ
xShuR6SfBg0ClFrwNMWmG9JkTV1WLTl9eAvAMq6VDXYivpKtr1Y/QPfYLzzsEsYM
gemsavHhTFJMTG87LhWQp+cKLXU/KdGpa6cazeCuY27KAFv15xEHK4T58zT4WQhh
PcDSnL0N3xqKWo2wBMnjHxZpt+m93oFk3fIMnvS4TYQRo+NkSK5LZ1hq+bK0kpSH
qwrRUHc/nHAe9VUHXErsIEE3Z0WCfCB10qJUwH70i7gDBzlFcPq5vqo53c2mjPWR
f4eRcq53FKf7xoZ/HuvirYyapDpth1mgWzR2X3bShhZVEQVtWJp7qQXNZhDw/7OG
G+F9Yx0gJwZrSHQHGYaWKfvmZZUFXVkjXSY4RAlASKvqqSc+hN4T/KUugdivti6U
+MpbFbpjtVYMfpWf0lM6IZCDlmcWOyoRjJKSRllMu5eW5OdyASXSqFhieF9vz3ew
tkmFH8EDB0M6bYL5tOwD+tjw35NYzNtnM1MTNvxpQTrrcKP3EcdD1O+ekHrneNvl
2PF73w9smR5hbaj7Sxkha3KfZE0h5HlKC2ty3+JZDbXAekdivco2BHSKAyB4HBtV
jwdmXdEK7JgFUngfA6VUoagIewtjiE4yrm69b3Y23GN38nfWLdNaztCM1I65cE2H
i3740uqa1Snpu8yFEspaQ1JfqW7lx8x0KqKTaVoGXGyZ9iKQAJeerfxC4ZIx04Vr
7bu9N9VTryt6LRP7KPH+LpCeRLGiBl8DSC5/kYHc2FA4tce2IJ5Qkbp2ZBM7BqT9
4GfezNOwJ3LapLrdlnnTrW6dXeq7Alg8LmtA9cK/5I446ctBsWEmQE+V6ia7U+s0
J8DXEI99gYtm8TKXkYYaZbyJX0U7570PXbOLFaIOKu/5BsLx6MmC7CICD0855t9D
ffmVF9nx9JvQnoZH7XB+PnaBlXtp04mpq01MDMy8fpn/yb3Q5PHYRNemieSpCLnV
xwNiJCdI1VfpUFPiXqLOruAce5S0hgtQBwYGAWe9qwxJaUJYC746f7V2UAeiU6Tg
0+1DqvD6YIvaRzz9b4GiaVH7+eqlyY82/jfLWDNtT0RhkdcqPvSC4VmErOZBneip
jzRZFiXDMQqEwLdoZNvur4jXN1EmFG4kSHsiX+SUHeFyIS4wBFyFZYw9iI79VGAo
cgWgO9DXi4+eNDyB/wpBTM99f9bRKT/DVG9ePfLEfDhiJBKzPTQF5qvzl3BL/JO1
sfsGMicfJP3xs8SDbgwiuze9wiwXP0Ah0z+mKDIyfBQzNE5tSGmlr40ZNGI1RtY2
f1A9uX1ADZ1r4Bt16ownrU5XYioVhOF9yxHFtA6ZCm2yW88JvLHJkQkSyq8zEyt2
LD0oSFN2Yq0gF1FTL/1YycCvj5Kxe1DoSKLEQ2dtjCJjQF/MShYe4+oFskyKCLVa
jEcijD1UIDY7weT3gMxtQyoaeCIaq6VjyfB9TGj4b1xpEtdv486+L7d5C+mc9abK
OHHbdDaVbmj/qnk/fhfBEUdPBONJy5Q8iYgT4jXqiRKL2yanzCf+S5HvmvF11Arc
J4nGi7PZUy+RyFj5e5VYk6XEvxfJ5j5fzuQ9On58wAnUOuwrwNWTkNSRWQPH+KdG
JF1E3LzPy9a9wflSVPY3QkTe2f5ZNvSZZ6ncbCg1CDsehchMPQhXhPKyQMrTnAJL
uiona7/dMwcJXEe3JBM3iAsHn4zs6tPTP56koVXOfw8B6lqSBt7tTP2VRInion91
r8jhYPoWA0b/zuYGwQjMPseJwOWWL1YeEWnBBmQakLlP3EaCMcacFw5IgwxsWIjZ
F9e1CqH6Y24YD5gbAAFTij3s+V1NxyA7poUObLVBYI5c//Yj998zYhKpZZgaTsL+
KceEn4GFYmHeOhpwn5elAWQQAuM+OU16Vz21tv2Vrz9adO83cUySClqKsOWxVY7+
0f/1JEzwmEHolQjC3srOlp+C0QgSef8iAf1TfmF/2clIZugyey7L4F260uFM0Vqo
uni3qi37KTVv6m4ylZBJIhM393SNlwh9KzgwVPIhmQ05LEGd8EkWDOdmjBa1Iu5G
OV9F8jwivUUWXcWifWdInZneUbhUZ4xZsUvSlzijrlzpmRlUYrR0jw0GXWU8MGe/
y0D9eHyRnNbWpwEjsTTK1mqpw6Plx1EC+Y7+J8b56w6JAHZspUi869QiqUrOofP2
g1wvay1vcwGDHSvV8FUeJw33CvSuDcNWM1YhfDDPVvgQ6/V3Z1AwgRRkwJ5l9zcx
0F3++b+1eB8xRAnEUNjsoOQwestnABuSZ8vTxTktru/kYjxLioJv2av0ljLqLkHC
bOH0ExZNodFVrvm98N4QSqIpTfDuq5PuIps0RTIBVC+unOyLwT27Va2niE4+tXLy
AX19Cqma1qFYZm3qiIt0Hwy5/OGVG6hnwlelm2OjjdmTR8XYyGtEa39HoWXMZo+L
hWj3d57DU/qeaIjl8TGaR6SCbJORsL8kVK3bX1YhaCSfPA/WE1gCKBRsPhQwKTgE
1Uxm6P+P/BJaXzdzhMLP1G5wJmpPRXgn20LYYfzqE1NBYHcn3seGV75u39X/sTj7
tiD3LLVghoYq7C6cdKibYPsnG/MHyGkFlVdXm+GcJ42nYQKTXtYbmHrrrV0L8TJZ
j9STxpPkSIiTEhWyVBquVWoPIBeLcwzJnbzQyewmA/NxCWbsCsEI8AIGdxWD85RB
kRQHAa8qvBv+gcEQW/yD4ViX9ZbFQuVExrCGtAQ9icwezMaYefVTAaCJWL121lcX
Ct+PFDUh1zHzoXMqDMOAktfRGAHlTYXxAu/v+wHDdcKHt6s7S25WXGB6K7rXY5GH
4TEPO/E5MQGLYvyGqPUNL0Zkbz0vxgeHXEzJ6emEl++0hHr1aX0wc+Z4QhZ4KaQc
lWTLOcqNEZoVaD7et0iCCq+eFwhniW7rI4PWaQcX8A4TEsMNRDqj1NoTpRwGM3wX
lSjYCCpS2UEPjp9d2JNW3uAueDEeR2gjPA7SQkLFy0VxxXExZV7PrBEDpN3LKne5
wJzBNpWXAYFiAQ+L4TWLtadl4QsyZ9BWu03wu7SOjQzCQlICSENzx87ieDUQaicr
14n4uGHrgz7M2602Flwfa3DXYgPxLmUjpJbkHmImcTcUcj+hpDD87maYSSAR2qXh
7tJfBfwCs8e/mCgNHPAC+BN1nxVI/YfAueIkhSnEDLp+ZVjagvH/xMemHx6ei8K6
Y2Wj8W2ZXJAIoq4lrpwSlZjWPBN1zRu/jVG/Nge7CrC/1I78RdS4vjsoDSp+B8ZH
kM2W45Kjj9kl4GOOa9O8EzheLJLKiE3cI+iaK3NG00tpC7wkqd2gluWWGF5I0V4h
FQNdq52Mjhk4+A7Mx+cxYn8HQ5VNsOC+KoLEEYMVgo6NlMjFM3g7qu+DjsLeeMFL
CTklHOG/p6uRhzb49EAg75/rBeUsF1VJuajjJo9S/Gq0VmmK+nE4654RweNYh6Q9
zf3Z0ub//Fkhy3M0YbFr0fjzfUadJDnHG4tVD+aWsyIua/KkfoEAKiC0HKYimq3P
8MC9HoVElJKiN6aq26Z+Py20GhFfcy5jBCbo4QGeT8PU4MKQ/oIJrAW0GUDbsllD
oF52Rb4V6cgnOfTukkOa7PQysso11JGVqffalKt2iJdQfCUp5QSOhsi0BT3zjxjg
VvNEOv6vKAasoPr9EwYW+kNrsN/4qybCaQIGPBKafgmZdjPqdBG7E6uMl1luE3bN
tNRgGwj4c2F9nIG5PY3uRYEhIZ/98gDg1pOAAB/iQxoi2TwLq+loxy4wvBnDMQUK
f252hdugFafSZgx+O/lWB99fAjkmuER4otOn4uIHDju8GFt6uExF85QTKkF2QU6W
qyZ08d6a94QsComem44O78M6sw4XIi50XdZIAVFTGMWTzjZy64Lc57uYV4c8fQ2x
Jp+uZ/XutChsGmTpJ3+krWHWw09nHT29iElMULBZ5TyjiMCTLHONHPLX82aW90Rv
5xjGLuUKPuwZQqcvZflFCyfQirNexQNeT+1U1JjpGGsWn99yMKcHSsAoXozNNync
QgEDpiABfG2zb1mIpf21ysWS1OwKb2HMYkGSH0iXMF6lh5FPsmuPg8ZO0+57egfJ
MXgvxZKiTBWCkTa30ogsGZVkriCB3Q6We025MBEf8T8UrLgFuaqRNnxARhZou83N
Nq4RKb/522FqRrdJSyvSFElGCfB+cxw50Iw98zVfdKVb4/rfYZ+b/88C9HHowwR2
tXnHBtaMI6V1v1imMZk6nIPAZqAId6IkXD053OCvAt+5PZUZlWkFHXsFSCSZZ7VM
ElguwCY0iZPW51aP9h6UJVuEJR0YBeLfS9QqmUuJMbbT2lUG4YoF96nL6PbjLxxj
1SPDS6syE51tQBAnkTI6223q8ZKR8eh7QeZnCwxbWmauzKj1gJw2f26EK14wuBnG
Ty8q8ixHNu2ONbhCQQAJ8irlH5HNrfMZe3Xu0Km6eo3+77gNn/T5N/53nStXcSOJ
hPaps/OUhSqgdEzm6M5S36b/CieLQjDRfFx1Gg21RNuZ4iZ6a9YnY409jlGBqtxq
SuAaUShKx3gTT7qvY9AQvpj4B8erzt2v2/5KwvFfZxfBixoH5rSWjWibo6u5N6Oo
FiHqMj/pHsI+IuoZZHt7VNbaibWlxn7/95XyasNisAaP29Ddp7pNyI+hVRRRxX3w
zNh/xMnFAA6cm1XZqZRgqWsBGNPgk4G0JhCpb69iJR6z/xpoIKcy3lwu26fvKfSD
RES+IM4EwVzut/qMpXU59SnVk5twib3aaxLhZwsbNKKMB5F7kxTi1oIH6KNJJqkl
iecDs5etnlTc6spci9mOZ+ECGImkdEd2SkWu7QzEdKbj7sZqAfiCGHVWH+IB9yy/
IWl3wZUX5ymtrU1JIR/xEDQWTs+Bgx9OhdimG3gvqJgoFVpBd63uohjskdxbMAij
W0NdHLlaJn5OkqJpFTsYBtSqUDR3HVkg4xd0yoq/okZrkRZ5+8GvEviPEvoS20bD
mLMiAm+OIF0XTZUajbP512lfLRMFko5/8ZsW1TrCcmtQSpGpJexkv8htmyBX9bBk
hGf5ufUxCGL76sRFha3gg95Q7DBUZRijK1x6Eyn3DE8P4GiLr/ozR+fZZ+5dr3uf
nCQGoB1mr5U/sotBoHSTIevv+x5VEopBp5AOzx8v4PrXDqA20RBZ7Z6NGTbR6B+l
e3/s1tiXxCx1TogWR37XBUUJ7MwS81+FmvcT/8zaIrFQ3fsm2YKI7H7Zy15hixdJ
62BgTUucvMs2BMKIKpVuESftntpYypm+/nlRtfJw5kGLv/UHbij/VfwVmYovx7Ri
G9shohXTANNfZsOwIEsCoXVaYtllMjUPoOabuzMkEyQT+8nVkZGzycksvoWTHUl5
gmi+RdaZxhzGxzGcyAgwIe37IHd8T6eEqqKGx+cpoF2T67VDNOhnGSUuaSJMNUnT
Zse67UndVP0wrhvp4wV9SNa8dnQSAYZc0HJ0Qg3FTwOBDltcgY0tgVqx1j+qat1Q
jz//GXP1WPzCQcAlsTuYhxjOeUraKVXNjQVqpr4IHgqJhG85qpnsj3CAo4Yni1Vl
jjjBYPEnWnc39x19AXcxcobRQQHmmCkx/BUBxH9IaUyodm+16N1+AFX5NRmWgi77
4E3k/sx3R40mymz7V3DEdaNMil5UsDwzltq2JwG8pvHlC0qdXqTt8CrjfPFBmKwy
g7bhVF8vtZjABIF1STISL0Ha3ISaCCjq2hJc4fGH1NnGGZCS3uuO5TMAONqG6RXp
3DJi/buoW1fMQAmVZKi58YAk7Y1nTnUDQSnDlMkcW8Lb3fC2NNpRyT7oXZtJu2k1
QmbblrsGBnwYnBtZ4b+Q8jpIYTdaOFIZjRftqtXHVqUB8+wZeaNRZLGgewt5uMwJ
43VO2OzlaMsUYKDs50bEuWElbOkfoY03atxjEC4lQVgvozmJWegpTQ2vEMXgjYHD
dLu5V92/VAOMM6VpYg1UQt1tMAqoaSCLXDCyLtbk9sKmgEzsIv875xZAh4tJkiYu
BOYK/QNU5KkcJgz/PCMnHnwej/SodKIRCDKgieZh/yuY58ckTrZoJosCUH8fwpoP
6r7UqitwuJAMalaxUJ7vSoghEWImcs8bJpQHdt5mTMBEpdI4NvP1WtTw04nFhl4v
oPMpbF1LnTBNv+E/p4HtEvkPgAne0MizbX+OwK3sUx1nYmEljBfozSh+Olkoob+n
VejUzAExAV2qXO8z1/va6fmtLJHv4mIAHNyiLGo9EaQ8EQTF9K1M0qVmmpWBYm5e
HXKAX4Vt4wNGcdfD5BajEd/rQlSv5aXwqTstShHDwap1sRBfI2gjpQCYQF21/jtE
/YF79csxJVZM8GAKyFGiEzhBr3kcIIPJ7u/Uu8CV91mRfrCHwgXGyi3n0YfE9ibr
OnS+CbdIorTi1yaeRFgAD0yhMEEeFRDDXf4oMzJIps5k1UId5E3nqOpKIPtwFc3/
GlnkCpCvsLIoDSNWvzj2W2lQMvOKovcdESNGkdaWfvzvL4Php3mtUawId1zz92ym
qCr9p0qPLdZir2fb8jwkBCLYmry/5uQ1GCZLrdQgEWVkJay1O9EwA/3AnMOCdtCI
+8oFcXHNWcHT9IX3tVq5mnZvzS2sqmL/W7wEkNDD15TCOO+jqtRxuiiKqpJd6G0q
YiSJyhdI7Q6+9FrLSCkQ2qOfJAfHHe4dwA1NBUg0gFnPdcBBF8eYu6TOReT2znJ+
CczCejcQg0y+087LdJbi/1FPAGr+aPsajomMOT9Kw4rO8hkVBLz1wNcgLfQ0+AzP
/wrP6Ey2q41vCofqkMzOnn6pRepil33OtUJDLzzKmYyLQfLkoAsaChHVSxMNN/1x
s92FrCM+5+GNKE4M9+pb+ZrkGu6pF5n2HmOyKsilpuVXzfyESzLKFaoHkk4swg6A
WE6JYS/ImhaATN7nAz1HpHgaSPEakeGLhdPTUSB1EF/SQGfuqFDViOhQZkPzXaId
uHivobk0V1qEKvEqjLA0AEJd6mGBv6dKxH3KF4TwRYqfVCQFECRtMTE+5MRnlskE
NBIe11ivhJX/OZ5/ONL/dSsJd8to2ksrWjV4818dFJaqsckfcappMZFzIIQ4qM0o
Pn9k3VyFYDKDL457ukyVGTrjfck8wrKlMwruZoVonwCw5dEzGEZmDCJZLnhaqXSO
m7eD3XnutwowDWYORTDerDhOAypcop2vtZw+wcZ7xSvJ1GE3iTlQu+cHh5+zx16N
PJ4YnAby+/eZvuOgEXWnHmKJ6yp9WumgFOhP/f/klAz6KK8j+b6axEdn8SxCMB4j
iCjtthUCdsyX7rktsCXEePAl9JzINKb7pIyNkG8yvqEVlpA6LSMhqi8xuJ0SBML8
MiPoPnbfkv2Ch/Mc0gvZO+9jNde2jumlNaZuWoFD4ocmYXWe4d60mANTPDfNrzwF
93kgtxPn7NvHhrIj3jcx9fW32AA28jQLBB1v4XO7znkPHtOgdZWrVCiYBO2mJr7p
V1pjbLgnLAoRjyk3V0KvuytH7DEMtum3IN+XR2aipBrqx5bAVKAjF9XG0IduDAe0
gbMJ18oXKs12X1n2BGwtjGqOjygRN7BUTaDdRte/eAC869EefJwNm25xNdAaMkcP
Ee1DbP6yasI47L13qVJ79CPm0nvEVch6edythctaKTbSCAU0NtteY1x3RNdCyHdL
79Uk47dCMejU/1KTsHKNZrppcuEkMTyS+IfaSuurNfSNMT5Dd/5VNbiyTVPLWQGK
2I6tm13BUlqENfirOYb8GfHbrFREJp8IE/xjW5ZIC80dvcEdrR4DFpjv23VFPwPA
6n704yN/EyFpmHSTEo4tvgxwSEJLjgGsbqbWVVM0DftF5kYSco5Ceyqytak/d6Ky
tvuVaU1yPLVtjA9lWh/Ron62Oj2wEdxmrVa6B6JRI/Ibu+RKh1GbpxRsux8cW132
2DRljqExRQakxPTi1XzEfxxcOMrqHMMybOCvC6fBFTG4Ei454PbRLikMDbl2gVRw
dH8KcdWq6U5pG+HS+442NgvGeFQ2Tn/+xWl85imaeoyRG4RHp2wEi5YyQK8MaR49
2TI+w4CLzYsZ+uuXrDMGNLlLPrtynGisp1WI5c6NQAIBTumDyAmyncWjfmcTrAxw
+STdm0HUw/WRHNIPC2nVZxroQfYUCGvzxHdmj9mT3vVHK6XlpE+MT7DmF4ZmJETc
BEi0N3cx2p2lqY3PTW/tOAG+1jyhrT0syfMqFxAveMz/qrU8ajV9BEPvYbiWmj2/
8/iymVydzfabptNKzIkNv+De7cwmRt4t43gDfCyy1Df0RozymI56jHvfi5ggxMfk
qtQzZcIFyK4pzRCaLXhe3l7wLsuHDJvsUFS46fktyhfOeRpGIRar2anvyZTrQ/Qj
UWDzR6Wd+gpJ+pDpMoY+q+SNwr/DT4u4D4fIsYDCs8vsYFphAGIqOM4vQi9zcgkr
b+8dcaVhFZRcoiW2aAO2XFuZcoDpaQIDOObO9MAg60JvD1X/bpT1vD34K5mKGKrT
eMEDj6aHZ4YU64DvBdL8IzalvCrLzE74bPYKXjnd4JeCQnzssr9YXdBaDOZFNeYR
6rUdtmPNL5oIO3zlS845TNLBTMPlULbaH3d1ihYAUbnmxvNu86F/i8HdaI3l3Q4X
kVdiqYpvnnXoI7a0Ol0zpcp3lp2JDRi5IqN5SUbi81omyFP1wTj25MwLrPvPMagb
IomZvaMkx0dN+B9tcrE4+c9/skvZXmlNAJrA2h4KnfFVhXhFTuyn4jUNBaT5QBTw
+oUEIOJ9KwlL6ZqujTFhM01JPapW1wFqFJpEvxQS+uL6mSWDR04VNOM8i1u04owL
1Z+iLntP4/KHJ8+M4LYw9QK940CHwYH87rpkgm5yeD3mkE7jzFcuwBEZpI/WCsEY
m915IYSklOGkn/4D9LLtS39pg0yCxBtQLTU1qUS54a8Pg3Rb+7K9xcWqTsCgow7B
WkNA4c1VKOUVsule0amikjAu5NQyua3cJbdrB8BD14bWCEUUW2msNMQInyNAZwLX
y+IQeCu8BE1WnHG30kguMUPZm/CEh3aa7ZkZ361xlowWYlCyFLwV9oSfqUWnn1Ze
JeLZF15MpKnicilJxs2ptOZqK0cCeTgA4PZZOTNbhT8pAvJZWh2Qc9LGZrHgmlfb
pwgXmITlFOSNxqPorpjq0SIeCGMoh4qwto6SsCC9StxUUpQstUZq1//btqscmd9j
aCRFsCFKWeff9OSH/osxZnZCp1tJCv3ykGq3SLsAWgvu3C/agHLH5XGTcyX3dkwG
vRxGEk8j6g44VEOuSQdZ0XN8fA+sjpvOrqztoBYktV6Nj3sSXCWkoBzuuOVksE+5
Yp9JTHgZZa1JsJBQypVJOC/nTEMExbeyjmpoVBaPCwCrsRyzOt3LyQs0pmmWNYes
FBl7S8d35eWUf9R7H8rbrpOnIZco3iayxkoJfzfykLztV8TzQ8Uh7jtW8dNj4q0v
vtgqNvxiUJJfoI2orwSq7DtQtdBRdGmSfq2H1QGozEXIvJ174zgPehkSCGV3TpdL
2RmkrXhSIaoTBUmGePidDUZ0JYyaeb3kxXnw74s4SrtsSialDZjdR3QEbskrY4+v
H1/pixY4u6R0QfHlZOmHaEcx5h4iAv02irMBDnoF/pwC1itf4QXIUUyPcGKQ/5Zp
MO6v4j6bQW4DNfGE09Dhl+3vGaK/7XPXW8HJgCTBmSWJ/WG7Fi/xPsNHCAFAgacd
QjsGnT1PW/2AUPGlsoa+iCHR+tbj8TDMGEAUH+0ri1iEqOhD5Ne2pxI5P32wVKFW
1QegvStgwX6W566Q85ByROKqZ69Je5BIukKssL4ZNrrztQwfJ3Cx+qJwPMQJe/KU
pu4WvoKOpc5xo/lphqjs+trETQ4ruZCjZLlfR14lsu/n63iavrC/Il7yFDkpfG/r
xgkwAtVoVvm0Qw+KCmxaUV6x4MX5iHPpy/4jBW1dVR0v2TGuXwM7ixSV4RaqTLk8
y0uprMrASnC0iZCIP5B6Colf0oQu+ECD9zdNjZACtzO6mMCvCu0bNrBDrPmnwZdn
vxUWTl7tzd3bKzpI3118sz3j1aIow8cu2IURuyBsEp9DrNB40/+LCqAm95ZBc17f
aSUHQ3KU2ANoo9v4VQxFHJb6HC3UW86m+xATIMKpx+HKTb8xIyu7TmCdazmmB9S2
iy3MYYdTW444osXhQJwkaQvvCWOF5LLRyq8NDV6S5klCbNzDdURaYFXaVctJWqrG
+0/OgCZjVVuZSSO/DOvk1BGUHiZFBLekMjpBSuc6sPzxpcDFf8Xx0pe+uynRwdmg
5HrMW8/P3wVuQfWPSa9Jf1HT3dqEVBwgOnX1w4dXNNuLbNXYGWC7anXrA38s2+Gw
1ZSowAsC21tQazHgmh7rQ1TBRN3IWe/r3zWZR7Xza8Vebba5+L3AIobMHGZIV0Ig
ccUQXjZx9V+U4bAGhSdzwQswbvcu17db53X73bbfIDeoO8AIhqcY2LnWkTpT+YQz
PgkEIlLwnRk9h0wfF4PdsFwI3SvvY0rjD8ILqDdzy6WRFUhZj+VDNNrDuPiU5aO9
f7WzH5hJoabibyGhmZpLPvvdKJiHvdau73drQrIH+MQ+p07P0ea/XbLixlK8+Gsw
EhTu+vYGFSZyqcMEYNe7NfZQ7ExpD33jI80gU3h3zssueSac+gvbSlcAikRiNLWC
oYg0VqxEQxUGmXjknoieHaOvUR9RCuOkEu0J/xtxHEdeStKKrfP26G4H1lHKA60q
Dy6oTRxQtbnt6bHUlwq64sA2ugVKmIR49aPFz0fun5ru0oOOZYBELFVW4zRMDp7K
rUmb6vsEdfYY+FEIU1NcYgKqK+MZOS1CgxN4i0jOHs3xn0GtZwYSyhljT7o1/xm6
+0EOtbuAxu9RqsK7fX9mv54MzgCWu0ShdHiKCgAeWzxU8D5a9wFsmi+y/Vnnp6oE
3GY9AF7CKuIcOwKFfVnXe96DnAyUo4C1HH40d8g2PBoNsqAu4DeYMTwZd95qsey+
Fq32ZrDrcjPrPbVkbUGz6nn1n1t0N+pEONCbtzsnUqUjXauWU+bzKnObmQt644Ey
XDiTnL+DuyJ5Hx3ttDmuUBcqsZ3UyJEcrZifIXhA/inpljIDGnNFsaqpY4waTFsL
DblZ22jORz8sHawsRubLzeO41tbWPblLpfPneN5gGq/vEE7jjc0mepEy7ZHScUeN
WIKGoc5ZSDzpBcfOKm6ZXegA4MaWYY+caHu1vibZdUw6vL/7aN5LG+QwaGu43+M2
xu52KDVxT0635+I5WoWP2BIIjfmshO08laOsUs1iI38/ssgb1Wdm5Y4lY2MHt64u
8nko0cPa9sSBgmxSJYXB2/Gq/cwnCxt9iotGFGxwEKiAexPpGgszAFWL0NDooGUX
7d2fXZZ7EBLK36ktuk5leRemUbbxUDcnN0aWQ7Q6pz4r7hlMmKbMnVFGb3v8+Pjt
vpqp/IByQZmtpRMkhiKCcpdipN5JOAsNw2HUg0axJ5ZbyykQrmgo4ravfs1dlW1R
gsAngWDYMzR35oxCyvssYlThtdDfynK9KIumJSnjmNtGJ9IMaJS4RFWs0nK24WCu
wDj+hDbrxRod2kY4xnCBLaYueH2T4lUt+vF7qckuM+nuL/Px38PWcjAJLZORijTL
C11I/wuLF1Cm7rW+1PTkAEEwT+Cn0v4rXAhhr2N9UwJiriW8dkDzyuhuLUxHBrJr
EEavg5Nin8FgFeBqyuOwDmomtRdPadSSnCQr3KUs0IpSqDjRZe+27Xa9FNDYNK5G
xnHGLJHyaUYSRLC1G4747EXlMQNu2252k4tLvIfW6f2pFQ/mWTg41WzBYKwi3DBW
qYTxS7Y2DPCAtV0E2rNSjamt/H1crEdYDMosqVSqbYvshaLBC60R/kfQo4J8KOFe
zQh6BZMCs6q0gk05XNR3BGFpTiSutdt7DbA2RlPYG8fn8laQHhLS6BZrWei2/8Ys
9Ff1q3GM07uwq8K2B0OTCnarLnmdvlD6GZmhcDZUM/rlHHpH/60TjWL4NUu2wAY9
5TwMM+VAXEbZZtDPpcJwhcQNn3UsHo8ErUAEwx+u5wrTRYUj73s4wWTOfuckYH0k
N7xiN+Bv+I+oCdBh3BDr9zLY3kMnFuMtKtaCP7GzfkzlYhNdYye/muqn4G3nR3fh
KON6p/LR7fo3fECz8Pyy2t/NefYkpsLq2Xot3R5QQcxhi1+Pogzqfm6OyR+s3CkC
ON+TCfdAAcIn5TsCmlzI50dZHwZpOvzKX4LczLt6/EinIf1DafpptJ92+P3kidql
6g8T6SU5S1j62DoaqerciGyjyyM/eRsC4MbVj4lY92iDe3dIsurbBFRmWyt7mMGZ
u0O9TmtjoWn0ZACpv3d5k0LbL8pioWGUVdCZuAI/d8AX8tWe9R/CPvbtEQ93AMvW
8vLAmAoTValdiINFsw2GfRzGxakeTHl8QXwMP5FyF2uIeHqwQOuqHLRuouRXx1Xc
OZ5oga3pvJbp/GsrrmZC2IbfU9z+cEOYpOr7ver7hJoM2A5HWY3oUJ/kfz6+sgj/
7PNGHrKi+9mluAkPthxv479LbrPgOCtV0z8M4eGARSa4cEB0jqLfTqgTMZfhHPQY
wg8BByMgGkGH7g2S7F/AG2foe1l8GRIYY84sD63FkXv6kizLqDwZC827dphNwJ0d
0R5hDT3ZeRMmxHgWqw0nZ2g7evN6/YgT0GFNJsCSHkjRURzz7dT2kgubglue78GP
gZgs4Dv4uJD1ylXXOfbszgxjn7ZktJqndJlx3EbcG2EHHuVIsIZv4vOoGItznD2Z
vtRBITlY/lxPakN7PrViQODZxa//W7Yl8IPSc9su2ZR4+WAdWjNTK7CzjLAYI0Wf
PsU1S+i6wwPeCpT1rpX3hYAztDn6NO0eMbEDIsq5V4Jo69rQD9/7eX7QrQOfaKRH
iAc0SK1CFioPebtU+XtZix9SYy/JVxg1CPMKuFTJ+yjrjtO8C6Nm6MMc3TuHcq+I
yeJDBP2L+z7jQuqLCBpld63foCpNg4l2v5ZcObxXcX6zZysV5cnJsNSNuH28sora
gxkgnTyMo2PE40AeWgqxzw/2ZYtSJeGI4bWyeQO85Bnn4j/aDa2zBSgVan+gaCCi
1Npka2vNWewyAMrYOG4JmFXqhz6/kF2Tem4lX902ZH9vmQQcAdzekWdI/aC/Rcl7
NB4yTJl8kewo2SO1734tQ8NF4Ci0FnxX9KiUC7AK5s8kTrc71AZvnrKVMtHt7DpP
uVfnnUOQpZB3bD6rDi7xjLWY7L8GpTqOlSYvKSEHje6dbdufJDJjKhZPJB10K/Yq
n2A+u3Esaeh4LBVl+kLiOVnhKUny2xbl9dqxcZfsHv1ljRliq/M6DtzrCcdJRVCS
ewQzlT80MzUx0HiRYlu22Z6B1DJt66rFCNWUNXHKYbhsy83/hAlRRnoPg+jYdJpo
i9MfW+oHJwmyF+8/tQqrW2dVXSOwHtqQ66K08DSqv6z6Efpu4vA381GqAwK9q1mU
67Rd5btjI7wv0Qwj1zuJb9D6myHy6RhW6vk4KoC3MsaifDH6jT6Q7QSQJPYYsmPt
O8dAx8Cl1eGs/IAucKM/qnv+9Dvo7n9PYSYINPnA2zRwzoz7+PsxZHzeAlN8ropK
x+FBi9av5WW5lnmW/q4H9YoD1Vw6GWrTgptM6T2K7rNRyJ0s4IKsUNhmoYvsOCyp
0xiqfDfjOlIlgxL5eenCeKAAl/qz8fqlxveQeTdGAu0YPIV+ZkfeEGII1/GH10Ip
lZEfiuC2A0oedbDoqpJQ4dQ22+XT+E5aQSLD3R1TpLISVq8YebiQ3jlJE/2QEnmH
lnQ4pbnWTL/MIK4Vq22C1uBVwKBjqSguiq35CI466bYYK8+U6nQkyTCIR6ojRDdm
INPFVRDfYx+nYGoTqno7dwu1+vSrjpc5jXFFNBtcqOAMZzgxfUzSWr03fZ2M7Ode
CyPSybIY8YcHkc6tHwxZKDEvAOQbSZqaepIzH/79J1DXWfbwJ78vQfyWdb4NHAfw
17QeqspSx7j1ASrd8XVOA9+Iq/BQBYaLgC48v5odN8t1iOGx9oak7ZibUKDbq9DD
JsdGnqE7izgsF7oWMzNC0b0aMAVH44p9Mh8Evcy8ZEHidx4vjAtYc47FMdmb/DHF
EKWCYGgbrT0/AIoOjuRMYLA0O3v+Jjh+NVEBAUu6/YRQKh+S4FtNEE28Laj6Mx0n
k4I0X246YSnp4Qie1/WdRp2nswQJQ5yqIW2PDNklKxMqPXfwbMRVCun3NTThKsjn
hcyePrlP3HGXfJ62G2laAj+kMkIPfZ33Iv18/iS95uCrNSkL67ea7Laz/rpXUB72
C1U2ITZ5EpvhWe7oipUX5cQPtQ9GaNuxifbteRwwG8OfcfBDu+xBDAbu3IakN0Zf
FhUlCn8mXvmbbAq70Gtnzwz3bjKI0l58iftMoj0vOs4wYRhmABwEfJF7pdf/p1KU
1ruE4TOrLuWeLykq3ntEg+DdMdvEGhrnUnOGhH77r97KfCf1OlCv8w7c2hFY8rj1
RLR9niL+aH2TDT75N0ScaBXrjipqaiDXWViYTo0lkMODzIT58oKZ4qJKSMAJvxE0
6zBYwU+57a7+Jn4UqqkWFQbrz6j226Uqfud2bXMQNA5+qim53/Hgl5R4rPqInAsh
SrEAAinxNEoVqjgDt8vWB0wgaiJVd/gzbkdpSe5c4AnRFriIlZFrrKSXaHs4tQlM
w8pt0fIBx65Ez/AivB4SxIvs/Ij7neuwqvau7vwJY6OUEVRiQGtugpLu8EF3zORj
fSl49ctJshqCYf+4SBEzV0gs/eDtbEmGN7UDxbEjDUNn3r25+a1mg3QBl5iwuo9v
GRKxtpHi9p7jotzPSlPS3gaOCeNYyjk+1/SbcBWgj5w+1e4tkS9hu4V+MXorHcSa
7B8QWNbal+0oKmy8berQxNmOjuw/uikcIzsqneddAC/41nTj+5j8YmdnCfVaUcGK
MgjM/oqIex7DKCRDgccofNa5snJ2+W8ETt/NXi5ATf0eTn9B3oNpWXH1m8gzTMCk
E6LOwgxTt/OiQ/z63PpkObWiNdyMRhhIpQV/pUo1fI/+YEdy86qKYeKPsFoBlYb8
VlMbRfO3WonmsIG6i03ieoeThyB7hxqn7NK7ACuHr6D9OkFFQPrgy6h1j/25mxyC
WyDO3L4QTiu8f1uTaxgUfWzWF02qYCPs8JkofuQA3fyzsTkoqU0vpM1sJwIy6gPp
j5o874YR5uc5wVmRSgElm6Qypbd/cuwHXZGRH7ANmYHlvwz1Oun5rECWd8o4E2cF
0FbPYA+WamRfbQoHGFqVugVqNyxZgah+Y+cRaF26kg3RyQ5QKHLfrIVH29MvBo0q
/ad/f5osvmIwdNndLLM8vyp2dW+Mgm216PoaHnUsGaepI0Gq+Y74KdSc7+TaRX01
PgWAc8RbkIwgUP+yqpd5iMCueR8tjQlSv+7NXuVT1i4mIY1fJAxm1G8YSuWN8OJ1
8O0aaxVWVK5FIA2Og8Kkn2UDg5R9yOAl/uYk5mUJargA1zMd0nzfVPmo1W8VkNMy
fsX5DE5bOr67Io/WhUIMUOkfbAYmnRqqdofXnIwNWjyCI051gTulqc9taWLuP9xh
N3bNQCcNux4RkTxhGXH08/iQ+a5nYSxHFpHhS/nMoq8ZTTRxeOBAhNViwGVz7f8u
paSDW0gIKKcmvOCJnIGJiA9soI2YAoE78iIxacLHESItoM2Cc65xCNKM6eXJFmL5
2WoSaHo1FuUU9CEPc+XD72n78K1+nFY1E2vVRjaQ7GqZHODfSvuLqhTo86LeZjwn
a1rh3LQHgAHmPUBTMargCOE03kSioHYXqzaol5IOdNPwfpB9YMv3cRJZ0Ky98wYf
jGTXRqU3iCGuxjuurSWKjkHiKC0H+TCOwPbBtWdpNwHHB25xU+P5CFX0XQmmUiXX
1PhDF0iEAWxgXcu6+GucdkFyIsKZdB8FwqVaLOGLwyQUFrmo+Ou8ICUY4bm0+Xbp
plm9us2BIQzqtolY4enowfz+DmI6dY8OE+9osmg75FKTGr1PeLpBpoFQcJMduXRK
4/aNQrRlj7UwzNgrvGl3L5CiDvJxpwlXkGfrCPMD1OtJzRbXrn072+xXXun6u2ZL
xxV+GYN99hFcg3vKrUl9DCtWJtAd4HedEPbtKYRpDq5rs5Ij0RfSZuLLyXSAdHmn
jt5VuC7sSL+e7JOHXjpzno+HXQ+DUrqhrX0n0OqJZ+4qZrquULANIsOAthF+JlBy
al28kSGoUv+6CIaat9HvS33O7UVeLETF5wB4j7KtdSTXAVCUCd0eBq8STerAgraL
S4vaPw+F2VC4zGetbL0XFSl2J94qXJYNQbdy2eBlOYSrHyR/fIJXg4kpAgwzFSYj
7hkZwllEdobr2cklw6ryeGr99Mpn7MD19PTqCIFbxGu8QWIZXzzJ8KgBwZSh9E87
Q/p2Qv9HlCWsu434QbzkfxQR9kOqsUZMtdgkP4zuG/IoLNBnwQJuWJbqgmDDMrnh
SEi/bHueCTcblEboJUgHpRoZZpKjXKQjN1cFztwF1KDGGj9aofh3VJf5Uoft0Aq9
8+5nsCbGGXYnHbQyl8D6h0xx9yciZ992buf4/VplrxzHi4vcyxj5mfv1RaSyUeJc
ag4vQJmX+3jFiwh8b1GIKhSjEv+5Tp2V9eVMDxmeDaAXXzG4buOvWk4W6353k+TP
XzSUpnfjmE38kifjUYvrpA33nsz1iQpU82UpY9PSBtsmF0uEkl5IcUH/YUUyT64w
sjFAhOKbMAa1k0gjKmqAh7wSQ+Bf5DNHK7XiGQdySc4Zj+dEnwsY/3zsLrZ38osn
IuGRGPnXbsYgqsEbaZjtBOr8CYtKCRyPP8MBl/uN/TZdjYRfHsXQ3JeFjppGwDTA
p2zAmK83FEvECS/RVoTgE48rBXOQDlvQu2FtbMyIEBLYfRyBKClW8HUFFeluQJ38
NaLAqGKXIE7NH1gnZrc8V91Bl6VJSgUo5mlKwKHr0KmnNNGEUeVUXJLccLyeI5vU
Y0qJSGiUCGDI7RhbyHOa3kDvNpEJxYo6sXDN3A6UIU+dXdCIzj1rp9M6z5MPrZ1/
n/wfRAKF5t7A5zqy+pOqMQCDbjDUrGZACrkM9yOUG1SBzGNsWIhivnvHMef+EEbD
NrnkQptpf0kMxZe40Wo89FqpRZW9qCuXtk6GxtSJ+qJdtvyB/b5dq4KdQ4DzkoBc
/K91wauafmNYcyGKmSlH3l8R5NGOvLRwAX03EOUO5oPHkGgGF01+YhMCB3TFxDiy
iocG71l0b+hrNldKkAdfk80mwEFYE4XXQJJldPW5MmOYssfltXh4KoMEbxSUDuTu
WZ7vZsIKgVbLBTzksMBp5Jj3b8d+eXIuE2/sy2Ylyii6Y1v5YuKgXZ8nVxZ8t+g/
nKuZizehMqnbF5x2pAZxCFGkzUs5IpQkj0pPjTRW/buVXPXnhinq94dS0RIUc5Jk
a3oRVFW5ECGg9wLpBgfWBzYNvi9A2INpgymOAEQSPQ8Ro5YcCjNu4hr63nWS+S8+
vQmKXScFdJatQlljB1vpU/mv6a+VJy9A+2hoYakdt4E0exfbATltcXlS8k6YKq60
Oewu3DWqOHpzFeOgM4hZCF8winkDGIkqWw/ui/PCJXFBwILf0JFHFE7mYbhBzSfg
Bto0FLca7r/bDdQ+a8tQmE+be8m1zhamXyYTVyqu05aNp7CvL+Ob5d88eZvhFXfI
TJZINesYnjWdyf2Ck56ZFkGwUw2GFwKXuLVgBHv3LxGLR4L89jmUFNpOJ6JnucTW
QPcZYaEkgfP59I3drwvLnpm0+/wdy8TSyfV1UgdGru3SGfaCPovJPdRlVveZ7qgk
Z6c1u9IKnNy0qIZ0B3BDkmq/FTsR0IKoLVkRG6WFOw2rXkfHYmxX8MfgHQIligP6
sp4r8Eo7G12bV7gL1UEa7jbSi3d4hDRj4+ypzEsHnWxWBhCzV6zzQe06IR2jjzuU
LbT38hWuLouL+uQuJbcrsdidmL/pm+3p8Ew0ntHxaZQ4LzzRKOkPp0/um+4rIm/Z
Pw9bZcDqPfEfvF/52iu0xNSkq3LfqTcHRcGQsQV7JINZFaqXcRPi0UK/J06Gv2lK
8B59D5emX2wRaqVLwKvuVjpZfB9weqYudCTb1CGTcIx2fgJw0oGaPW40lAIBJfAN
BVDTK/Rk5kDJkILAi6v65v4S0ZSszj5Texw3Q6g8AvzLHnyuPk3/YiwyM7hJ1biM
517hXmd4anq2Qu2kOtmH0JCyINozvXBem3uGlhStTBc1cZCUYNAYQjen13ZkCBah
cO8PZZ9QLzaFaHMePfkY3wWoqjxQVoCdp4aaUfJR55KKsfs+W+0LZuaX2MkOyBKC
mP/xsBHZxUdumG92jHKpssK/eP5l3X8hnkFG29DXj+EU99qqAfEJpbfbUeJ4dNnS
ugOqlnROo+q4q8nsJe5OJapLBdRDRLon8LimxkwxHJhH0hg71HjhO49gB4vH0IK8
4MaS2xid/VtbCURoqkTUivqIAaHSNbW1Dod8SW0wF06eZ/zM8GkjMQRlrKFAiTaS
vN7vXnHeAiVLGnc89iJzRCKKQMXW+a/FCV/GeOxPC0zu2g+gJpEc9JkL5MMabhmD
8QHqL3pMQXEV2lRg8JXJuN0DORGl39QdKePclQqcXh/XM/4bzqWcTh2bQvM+IB1d
xfljjKBtj/4j6DycULAWXpwH0k05laAhBJDxomQuSGQdtsKcsWL/b7IaJ9ueCh3d
4wSui9FToJH9SkjyYdoX5tVcLGJ1vxF7ptaCXUmmxO3eXXay55+DKBULliS3KNwP
g1kpbrROij2T/xKdetww9SQ+ptsVqx2iVFi2IaUAx7NIGcQ3m+Ykx98ag+rk1Y1P
baxgAiBUzOO1RlT+NBylwHcq+dYbPc1oN0F3hctBQB3dKMrz+Xlxsk3Sa7vBD3Na
ODMNAXXvggW5N+mUgv2v90et2lYcGdQKmyZT3sX8KzSIo0OJC+QQGtVOynxRQLcq
q/Q/J5ZeP5OTFDcRmBp3NwOrlbwS8Lienkzx57VvjJv7KZeVCmIxSMwxv+gQJzOQ
Sq0WAeMYrulOv75+ZtVFZvzUSEqxJw8aY9MR6B82INqvU99y0i+32Va44JTfEVY/
hY0CqZ+4IlZ1bBD0OYCV30kASu8rvmFeGUyszRbuejm6uVJjqrSxMzG29lPX237z
VyaoQWerRyYNwp7i/ojMo0DaBsCnAXTZm9a7EPnlTn9rI49OOlQaUDxpjOnZKAxm
FycUmnVDlEP7EP3xxUPojPTX2SgeioocO4NZlvfP6klJldeEt0ngf4j+EINV1O1J
l/mGO4rPI2RYGf5DAQ6pWaIR2+6sTsl9Z5bKI4ZTTutNX1nHJflMz99Y9lFf43ZS
vTcWqHBbyHv+iPW1FslO2O91BR7L+RNaHDSVL7Q3w87xO18qsaLS9/2uS98MsN/H
BpGp6SNSYVQymLd2pOK5QHn2cCWqvPt2HXoU2cfNvz+pDPeH+J4xeO3hZgQutFsQ
UvU9ZhS6LoZs1B3TIXX/AQND9Sd2eKLm8b6T/FuBjqZeBuMDwKarRyNu3dsTtn5K
SD46X75MCzxnqIC363bE/keLoMLiOCR9j2E8R90RzdXGxcXgLbfKdsXvKY+RMaja
M6Quitv+mVet+HHXGcVtvOFqsFmzjIOLhL8jvmrgyXU05JqvDVC0BHdTqlmxgkPO
3cL1DSs2BOwiKaAAWbmxD+nbu0nUTNmqkJ+t3LvGUeCgx/O/r2PWeFp/RqSyV239
XrM6tSUXWQEUecV+S1yCLVfEyd+5PIh/1td5Tyz/re3458qiBTDJv0QmCfaj+WV/
zvU6ua5n4rRK4VL0XGEh6aFAWefAWRv8+e/xbgvAaGfTAth3/4XSd6EzlWe2qf49
JvhdVUOh9bxGneQedm1c0+d02Fjc4lyZMAutmjEynI+My82bmdYgfgLnB0CuDVUo
/6K53Eds+Vioy7//VcNpZqzRjlSUSb24ES4J03oDHEzk6kRpz9yfAQjBQ9gGH2IG
Itx7tPelRWHe9xD2esus9GCUP0lF8mWaIUXMPjrljt3giarhAkBSEv5/btzvzCWk
PeSzI/pk73ZsxVUUftMs2GGcEwnqLbtei3Ded+1ViBHOd4Rb8dpGWiIAt+XpOqQQ
+doIZ2HR4aIUJrumDer1LO35inKVyjzBFMZ5njyoQn/FnKCdTrN3C2DFL0L+m3hG
Lzm6bF2Tl3P9f++LcbV9owMI3+tLfDbT8p5BBBwms3znoUCFfHRabutOy7Yrz+tt
UZLsQX1vDj1twRXnRx6Hb/Il1hLah7moWupV3jFCqFctMFm8o5VVPNUceUJXz+lG
83ZSsHhYExVHCWDRwRWWy62Lex8wj8b12V72tKTjRC3aK+IyX0qyXxsWm8LpX6Ni
ZUbDjM+dpAtOSRITXlhtemSV4l8i1Xr1u9Guj5P5ueBL63FawJO+OQDvbPGtZ71m
v6wHKGiZ73E8kqwnErdWIdg6wIpwT9vSJS09oKsb1UIABLJ6l58FIJJf5CytTvbV
tw43QTUmNinQu+2/6/YbVLDi7vNYIr3keU1T7Cb3jSagQlM00RCKz0rkvTC8ZYvO
y57fyNHvQtTRTLZo2tc9mM/6WvlRuGY8ScVI4VSugXAtfC18JZLa/3PPriuK7dY/
xFtpsPW9sjTWPfu0gvHSaaapUSan2scoZTlCosxCsPnJb9/xeieIaXbh5V9Hn4bC
nL/F5acY8iHdRJElMbmpCTYXZcfKRnLBfo24lQS4FA5PReLwidSV7pG5ReAfJvDs
28VslNiZJX0w5Z3tNK4ZKhFAlb6kkqrGoiLqon0EWnEM/JrJbOsT0nuLxTO20Tv5
Q6ceuIJpqtrsg1YzwJw2YHmBiYHm+kmdTtDcD7eB9a1+BBnDTR7tFcYIp8F1if9n
74OfEP61JJvedS9cabcWe8O4WAtGIMqIpBCuXYnKMmRN3jerbKEKOhehzpwn63zh
j4poNqzvVh4ezzpTrM2MSrZwcwwKoLVbmNJxx+W/nrPTYRCLb7XZXdooTxYbKf9Y
3kBt1D66LXem8oYE3ecYcWvkHq5nmtb0QzhUy8dNeFEOftBeT/lnCe0KKMVew175
0u3hgt0bT4X8b6kKUMIdQV79rVnmIIdUqk7qwrQ1ud6RvyjFOFmkibUoQHV+NIH9
9Lzvw3zoHvfGES/CrwHkeUmlK6T/XSC7ZXwDEVHc/wJkFb0G78j7oeJ+6gdRDRSB
lQz2pTp8UfGtqyK/OE7chV6jPUJ7K2E3PKPxb1OSaTps8etzQq4LT7+407Mkzy7X
sISwmsmVff14O5RaInY/hc0mkmkYtsBhHg3zZPgDnB2UE2eXGZ+HyCdAgwX9ywzc
w48SjAapEdI3hZt9y9+Yiq2iiRK9o/x7yRhmWSyBp23Piq/Xlu4LyhJZ2HOs34wV
Sxae9XJObpArTNp6hPE+NYQEN+MVNAlega2dTQl0aKs0NaFv8rI+pNgM/zqWnN1a
jBG6k3nG2ymioH7BmvNHyXph/P7P0KV0iLTpEJDAMM23ovuI7yA1O7veMJ+cD9RT
Nwxd9mbtiQ829BkEgtWLVIA5NLMPnC1CTbxT5NAXiU41edN7intAcCadkAoLMxiX
6ndoo6udWWt+p3N8VyyTlEhfPGgpxqlqE1XzoRdjlRv+xOlROb+LRNDJ16Um3/R6
OBNmqzCAIguWXuRUgJOpb3M1plrajcHyULdsqmvbktUeQ8irL4gKBnZCpi+fDjGg
Xl2g+uYUATjYx+MkdCQSuXbvmgVnIYJShL3oNev/bBRdWIJ6nSUllGB90xvwDlm1
FCSl167hnVTmDUXTcrXwaKt7oIywlQ94dxqJnhs/BfDMeKYihFLw606GrLuaoGPI
NOb7STGnfUuamE/JXDj4tdNwoRWheQDKOk/BUSyfOqIDdesFPDFnOtWSwKTtN1Cg
HKw2efGZlASxLTy+1G9wjUhlPJlZUeyyK0agpxncLwzwLlS6fNQvW3gj8e3A7ilt
uCUXxhFe6rS5ncZJys/Tr1TOrkL7YF8CsicPbsEDHAFr0xHyJXkNylBOaWlCbUEB
8aEShCud796hE0rRtuxP8w+YBMnf+w2uO9JZwH+7ORkWx1p+B+jPBrTesuApwvqz
F5DBJWV9I403PXjmjkybAVbnoEoNdqEuTXlTgFRg6CjiDoLaZhvklDqYMqf8dkSg
7tCXmVuRN2VE+23f7DUI3F6QUDmqHdngToBWbSwxUY03UOv+i3UScJYZZ2CETPKA
oafQaKuuD/otf4d+HaHVBl9ypGpUr3dCT+Likey8VFsnYXytzs3Knk2YyGrZ8zlG
Cl3wRsH8nQumQGzI9YU7Z0iLsQPEP/DddjpF5FSKbw3Rtn35FjswjaixW03GRi2S
M1OVakdTp0cqnyEjnFJegkal7pkVzf+3UYX1CfTgBB79ITSfviVufPTCPq3mOFwR
9tmS4Nc7p18Su2zbvhDH8OxO1lB08fQm90kSHf0ixtXn2ngpmNosz3hhVQ+uBJ6c
+/kgxo3eISPyKbQlGxGTFLx8Bw00a9D5CGLSqh/Hagavtj2c0vxYKZVJ/o8dSw4d
nz9VwkWIVTnlrYIuvqkD62Yl5zw6Aeb801zCSZGf8zvltKoN8D+bDq5Fky5drtOC
E6XcgBhkX9s8SNfWYtCU8JX75cCkS6RSUb8fmglwUhmOiVd7/1qosrccuDVuLRnG
pcx5Lj2l4VAK0lB8CHxVBD7044Zg1yqw0Kfx3hmiZTC0yVfAxWx1wg/Odmkag27q
5AU/QkaJf6SSmDhJaSJJXMpay3h1rayFD3cdvShkpexFY9CgWFUds55Zf5v80Ggb
uGATjWCJOklxqnkHem3QBT65dlvqemUJOU4eorvG2pBrGEo9C3KjsTrUe1QKYUxm
4FX/4JXTei25ZGk0r91V2+n2jgSCBxRXBSv5AOhhoJIgwoiiQ6nUn/eVVl0nbYRm
h4ABATOs9L9m4s7kSoTyZrU4pFUKtb8zuIZqszBxj0WF4KtsE08L+wR8kPyTft5c
ZoYMHmXD9RJvWkW6TUEg079sb6NVMWM9CqV6ojMm+olp8PoTAGI9OxbzNfpiabY6
y55JBD13uCXsiA3ZMuAeeM7z7Bg4OJpz2bi/xAbDyX5oXzC0pnI9UrgFf3eNUobY
K6Qg0OpDNYwuCJmVC+X7E/d0MESuqXl0q6CqXWYl7Fv2WL5rQ5UT/ZPDvTZRi4P8
NSPJlssRsOXfD9JTsM+TD42b9UBAWqzsiot6FhomYzVLWdwdm/x0YtUltUdB7BXg
+d6PD9jRNGci0Z52Sl3MMS/HUzoq2nGBcioU0p5sqmsBzgqcHloiJ+gTzjNY2uYd
drra4wPYzFnriU6PoMZAG9J6MNS/EIaKq033FRs12LDihovkH3ijmYYEndNeBqua
DWtOhyKCQmauo3V9YqqbyhiCGL6r2DBuVK65fSkMQ1NUTBdekTyaYyI+OTlcKyAD
PJsqqVZIBQ4Xusvo4rXewc37LfdE0wzmnoti2d8mQEGNMieOczzKyTL9ZMftgiVG
0J3krJ0IvLk3Jzx2L0QzGsEUwJStq4zTkz9PwVoPsAq+LbM/vudzQei1Ldl0lObR
TOL+Cibh2nLKflvAMRVdYturxaSFdS279jCIhSxPiyCPxCOAkoO72JRNPyMupz/z
l2Y3UDZBo+s1fkSYUWCYDymJ5GKqMDLGnnLO1GlE68mkxAqnnFPUbG9hCFg12AEr
KcByf+OltkVgMjZj2RJiDcN/FxLF8gX6a9Jli0DO8434G+njfI+q9VWBpYzvo2d0
L1iNs6csmK0BFeN3MJow9szqIlI3auFgJq3a/23sswUv30Sbw07uJ/tvZpn3+PK0
SI5CFQgZwTjTk8gaOsNCXxXpCzxe5wNAVTOHTuXYPUElwfDuJ8s8Rj4pXI/3kKZQ
lEubWGYo71hHFJETiyGMstWNZcZ73OqfsEzjNjASofVp0Fx/4uc3Rf/dnzpuom/d
aae928Vs7CK/MmQ1UIt417fr27rNZy65rnaoCaSD3z1mBCWlhmJDAC6TV/N3W+ku
JHP7qdV84N7cpdUibSlO03pZws2Qp+fenesHqIsxTW3PIXzwP3RnGX5X7nz14Wu7
XrHF4JZVlq82YokLsnUsA7XSHMqaVYeYkzDYo/kaCFYMEjdQDvlO1/uyW1c3073l
DnmY8e1LLqkL1Z5C8Cx1yRiEBAcIIOTm84MEeiBa5cBE5y0mLb32WG0SILkIorGg
BvwdhJN641xWFOZMDXqgO3b9d7hnCabOnD/snMtowIKpbelEvqKUFTtuVVASChOy
iEu5HkXJFduaWXdx5widS2QFqIw9cvAmEy6Mldu4PhLoyQ51O3QfcFU0Fx12r0c/
7prqEideEvLpb4+uHqTtgTwws9Hy/Z+A9ritbpZxBpp1+ViJHWSz60Y5oz7G2Lth
dx4KUWZmRQ+X5W9MBcPoWfM6Ln14nJnk6UKKpAyLvxhqnZDCijSbz7l8qibq/hKk
brixj7csTE80duUm4rUZiA1gdksIPxqBN7rcG7y12x8YrkSFTH/IOY/hZTdW7B56
N2ITDHzY/OBZdij6yQm2Kzt+I6m9fK6l6lln247geFcGIcP58x05Fi+mjjxTRcHo
xECj0eu+8PEuOmMqaYxQ4Zj9Ks/stb6VuRlBCtUxqr/LY5QaeBPfDW6ptCVg6vBc
W5x6UWUbkkOTGEhyZ1OFRun/EMWBBmNThcmclFASvzNUZGDh7/xdyucqrDytZrps
PWxhfiFMozNGeY9srFr1PbO9a1uhhhq4eCFcuR9A7+rxHScRN5mKLRXNvXdesbkg
xuXD+2TTmWDYEb0ZE9faB5SRdsng54vSfSiAIUNgAkBAeZZSznj5OyvfFIm766Oq
kbDFobPIA4N/V2SATGcEp2mjXPFsF5JIE+A2JX7RGaCD4ccXDs2BeKXfLjUqxA16
grfekFYxXnBTSZD2k6FvGbbdkKhdJ/2xp7XxHyG1b2CF394tsG7CPLBFSAS/cw2W
KNvvoQwqssgoY3v0AuMWr1+awtsvv+p0m1DWxQQdmSsZpZYpo55+QpjOv/DNLrRn
SUi5NeWTEVgG5Oe4TVODWqYlMoN6JF4FSNUNF9HoXOi9G4QUSGDrwbfQ3eNRkonu
7rF3nLlt425gTUyt/Kn30cmBHVYdozsk7JN7lIT6jOLF6R3zE2Oq2C4ZKUPuryru
rL2pOkY13ZgrZNu7IwUgk3YomtwAn5osfqEo1pYpCdWf/sFgxVLognns1c+j3uBH
n4Xh7S6SC9wjoO/Hxm6O2rARRgWrqcNNHgUpwN8mdJd1sIEZHjZNhTdgIxdoXCeW
YI2RxnlNNSpmwGfp4hybyT+J3o6byY3aNHrePzCvOw7rmhnVXOxEOoFv+AJg3P9w
Qis1oG/MvXFqjvfJTKQgJ5EBoeCDcWf5i08YsMd+MU+FMAm8GUc2zclstxbkE5tp
TSXLU1EWmLU4MsWQGxBqF910jETfMubeRm8XQYub/lQFff/MRi7xydIb/nq+DDCr
m1DhHK7cPXMVinVfjwAygQ73JV5XeTh+CYu190cTDzMfATwr/Hdmgi/IN3LDGUgR
Cle78FRflu4ZSpprNnMTUtKXrjbB1KPG1iZ4IJDrBcw+F0Dg0oM0GmnUq9f5I+Yx
OOwgC3SIMG/fcjUrBVPlAOz4q+GxTRsAJ9eMFlxYD91LF/a4HGKPm/+kS2ciDmJ7
FO8fsxf13okdSioIPx8zlnVIBYxPnhf428sWhOeqovoiHATP+oWu8HSaCj710Muz
LQV5J8dw8egNM1hEsiwG0jDv6N/PlM3Z1sUGWa/9D+t9w5gKNj7FT1QciAACIwk9
wCOjQK6mLwly7erq35lkxX+mKk78ZpUne6Mu17PwCFxhMKgPDqJ9uQWL2MlULekm
WKi6d6le7Qv17ROypn/hNYa3E/Ntd7eJdyyfxgoOCyAd2Jy3MnFLE7a/dSkVV32J
58eTRZb9Mw+xe40RTefLOKEwOR2nb3oITH9O41/+3FNt1YBik5nbTw//Uv9et62W
lIHsfctUYQE143GcA7WnQcwz09yN1ADyCdmzhFS4K3+sDgV8T4MHwWcTWpXnfmWQ
RZvwk6lmWP+TIwCxwsFpl8sWfUbJ084Um/F1rLvBy4EGo7gyyiazifxhnrM0coMf
Yztm4D43UD0pCSR9DMvyDTShjKGXXhBvOqoQFaUcqw47kdcMMMJeXbBviXbNE9De
MnjyJ/AlOCJP9H3gS8lhmXqb7YOPzoXKxnWPK7QxG8fqZyv+CjGy9V0AeUr9GlLZ
/TiWbL2MyUiYQ4VfR4zfvWGndE/jEeGu3psyUFuu/5NlVisM399pYB+Cxq3zS5qd
WTPLEF0iBdOAivPwB96BCLBCgkqqPcNuQeUsZrspy0Fg29WsKFKmh0VG0ZogN13N
i0Sc+rabj4gzCvC27pWLR1llXZTSKXWYijG2ZvlO30Mh0+mCho4AkHRBln2JT344
wbhzImucqNFeEPT0s0HwQ2bfhpaV1hqaATfM6eTKGXtZ7zK/+YieTkoSGvlkcVH6
hOPc/vZzLW/mqWCjYtfN/mfrI///tQYhDbNKiV3c/hiE3DIFnow257as997iVHVd
zGle3SsnNo0YuUwHUHxw/vJq8vqGUCFyK7mPQYcnKEfb9UsaMcrPziyXj3A0UadH
GEj68HfwsXoOd3piyrTuqC23/iaMsFOhiuPffBBsIz/Z6hyPxgkyvwqBU1L6zDES
x9KkheJYJf6rsezgBByLR4gRueOw51mkvSb9JgCk5gvnuqZoqs9mVgQtd69i3cRe
Ylb1zYgB/BEkCHCSIm+N2zoliLzDWbN81gg1iCHUvhTnZQT9onTpv254joEOKbj8
M0OJ7tD/BSV/d5Ue/1YhjqE+kq3n5XqZnlfPRK7OBEwjofxQRgFLupPa4Mb+dRk0
IAIYBGsSy4b92A/knvJ6v+vLn/GQXGlaexAoQ+uwh9Wd0OgFPzcE3Hn57bz1Sgi5
w7dysBD34CyEgEsIbrZgAMLo+Tf0vG90H6rwNI3bMFdZbb2bRF/CVMP3clxvjPDJ
KfVeH3Py/mS/HfzlTXZV5u1XoZ66/+fYo62V2Ro0o4K9ZPIlJeFfCbSkfi57J8PD
nOCJk5Bs2IuqLj0jicYim9U3OYJ9W5j8GgnoVeU5XRRjkDL27eP5LN2nMEXQ+Pbp
jECAMZQAuJvedKjg5JRr9/jYVtIRCES601jAJNvXp1lPzgoTmQcm1xfh0Ey2nrrX
YlJra9HttsNeicyk09lduMMZupwaAZ0k1ob59+XC+uj7PFqtQEBNAVGVqxBL6WHG
uK/YKd58z7PJkfJlurzR35TPJ5J75Lr9wxzkH+XKb9wGzLBUPJ3892WgkuRoOsy5
Z5ek1up0hfX15hybuGuaBXt0wIGR7pDZ7uOW270yyeGStRsBjRGWtA4PxRS2jFCx
n/z9N+oEdL1/HUjSmx1+1P3P2Z0IEOkQhYutxI9zrIu8oVZosqYz3zUyG3s70MuC
sPiT9OjWZq8hgnR7b/nBqe8PvYPN9SkSzOv/208iY7KOsCPu+PSFXHmnpq3BrsYH
JNHQbMuE3zN2BEJMzfb2WW/1ESxp0RRAdRU93GRkVsale2oyGLEmo0N0zLnpMsSM
ZBKWsOkTY1H0tCsTcWRbkBfUCDclCzuJAVE32IPr3mS7G8rH/eKuny25VVymYaaF
TINOlBlwFl4hyV2Gjp/NAUtyRZOG+hyC4zezxxmR+WHv5x1qXb6fFUx4BVkcUoWK
dB03Gc0Rd1nJ+/12luEijvY86fM3yRLnWVUw8npkYmxKi+uK6XNTMNlKhAeVCwEK
gaCALOdnKTACTEcY6frUDUeFfGNFwyf9I90vl0v67cc8CZ+0NVfBKddsM9hBzrvZ
ppkqYD62Kio+6c41cnFNY8zQ39Ia8XwISw++dv/LLRvj+KOaHw86IW/PjFrPQd+p
lL2zBnARalLTeu+pJI9LoylXugE+MZU0ghidDhVh7gI/Yd88uW1w+zlL5CgJidvN
Y2IdGowJwgX8nxsnpuX9YwDu7E2db90iTE8J6Go04UO4LTYEbcP/bjRF+IKCL3ol
DtBl7Ojh398DCm0yx0PuV/xjggwSkdEGxonBCnSA4yLk38LWaRvtaQmZ/Prypuy0
EX9f/cqGOr7WYftMpeguavny2Rt+1Q/FOGAQcLB6kBkqFazkOP1+GNaFH8G4G8lR
XckLbBK0t/YSem8wnCOW5kMgqCpBDhj+DHoxKEYJTxs1HRV2+LQ4CNVYqGWTgJn+
jQshRfEKo5zIs9YaSq4XEazDYfIrB22x4TaGME9s9SAWY07Dci4dmn6iN9+mQgNg
lj4XfTzzEVFGoEXucGx/h7b3SQMQxM4zxxNf1BCz4DDy8ZENsg7oHj/ABESuMpJ/
1hWOEuxFYgbRIIhzEkXWdcwoHdvUIKQHkj13v+/lsSAbwjFbrNWrFKzAcgdrzEud
IjsYcClDtudZyOdNJlhmde7Iptbh0F1y+3YUXd6TzMahReg4xH3P+qgPS+PW7/ZZ
FnLMQDgcc6Tp8PguNYmXmWK21YdI6BTGfttzq4DdpCnZA/PMFJX5zto0GXP3KUDD
1GAfgfVPWmbVBoDRktbRRlWJcTpBO62kKv0u0TQbgmN/B6qB5pIhB6sHHNSOZ4uM
UaIHKMVyKiUWxJjIAF0ZTtgpH9dGSGX/0Dqecdr4PeaKjRL9u7yZ1bzJL35vqvYc
5/R1jbTAp76NKAE5eiZp6vRLL0ZP6Omh5O4mvVYAUk6r9p2ZmWUTRUPY3WTinkMj
L6PdwBWCYeviLQZnkAu08YA/q6TjQcWJvINXvG+CHNUFakfePOpXjiZXwVNYC3XY
K9PqGQ/Rq7N62cvqVYEyEUXHFtLTlonac066ZpzyDe/GcxoVMu4kYFdK5cf2ABP0
fdiy7PdOkLeEU58yH+7pKHsJKfVFFEnzSUrZs06kJLZhqgCevAHT8yFxL1fXtxFy
8hAulvpF1aBAHJjUxH8qX8ZF4jU7FExY87M1BZUIZDrLc0qoD+VNROYpYtieUlf7
PPZBLxljA/3HQP0xJYn2T6E3ZoElWTKQ4RcWcqeMywEQQ/0i+vqgtIticiBfDKTN
Acf7WnyjZ7quy3fF8PwDFfbyjETf/3Ik6CIipcy1vgsWeLN62rAw3IRGFz/NVyNQ
okg8MXbvkAGW5su9dUOC4kSvWE7oS4Jx7kwLYjEwBAQagM3KsFDa18b0qORXbsyc
JcFFvorcH1Eg94OVw7bsT8HKbhpr29v2wKZCG463T4e0A2bcaMyOFBm+J9NDdnUb
dSxZ2VEgYX7KBKjD66UtT4IpruERKIjVhcX9j36oyiQxXudkxkP6AOehm97yNRWb
bWABdCKu4eZPReFZ7i5qSsLgYXndSSulO4MoLy7GPjs/R+pq+oXWIb3eKdketxFV
6ySyF4Z313m5s7+6PE7wgQLOxgjpYLkllwbVL5wBqrGmO1q2zKHF9Z2YJxyJeum3
TXfBGGXbKfgOwdq0WmV0MeweYWEGOH4oO2QfOY2V3LNmuyPZlFnw/qlZ5erg/0h9
Urb6cCJO6dqcRd+0NQsHMnl6JDqio0ZW4MOBh7fN75o/Ed3BrtHODigJKpIeC3oI
utp9MSrSFZFKt3LLEeN8L1Um6CxbZg07VQpaj8QsY+MA3HPZN+JppMTxIGORUNns
wY40L+9OBxad6RtfHhmntHHZdpdpCPKFjrWkA7tEf8+zqx6akf6E6mAvq8SQpAIU
FBsNN82Uq3nTu0q/wV6wVQpBgd0KsoFHcJ5FrZJqH2YA/SbbtEF/TuuaC0gyo1Pv
GT7E+smRldCOZbQSNAIo2YVA3pL+a61YhRLjw4RMtRnsrrFQDcgZAYd10ATyUIoH
Nbv1YzdlIXm7SEWw15W5Dk/vRGNVdQOcn5p53QY8MvfL2SYDT7aY3irHj9X0PCIz
AdrwuGxIo0ZcMGyMnDtLXxSmpf+UMRC7Zw9QLi85s/rbiNLg1sdVhG+/FnDmVT6P
BsiKzrWiXqLZddFPYT9x1L4pqF+9S8oCkc07zoAta7PtXqw140TjKvqKH3dKig4N
0e0oYs7SSRxKWwi9u9pblDREkMvnGxScoCxO8igW4/Gihy5fMDDF+Z4PC9F9uZNg
yFTcYgZ+Evae9eo95Hh5Mfas4NLQPr3Q9m2mt0BjZD23cko4uvmDxqp8TkFUoruH
6M4h5puKDsUqr/1fF6HxY3dUZSBONQmQ6RFXom2G07A1cC5wkshB+/BM56qw2SUY
uvD8eM6BV9A0SZv3Az3JGaJ4uPcQ8V5lAHZcqs41dwashH/HZW+X+SuMBM9lIgl0
nqHkie+fqpu33p2tUjcPVWks3yWW0pAA66dX/mdrQtc6L3/bB9cH3zK3Wuj6TEy9
RXZmK0RHIr+LGEnBep1850sZODcteBR8weXMjPMaRe4wzrKH8tk2H9NWkhWHPOYp
0m/h44gYYgGNXpOHtdQE4coTdZTmT+6lLI92acTXx8FrY3JubJI/HSxAN33Lfg/c
5twpAcCc+Y/kO9FM32tS+Z7WyikMRsA/tRjHu3q3vZ654dXrValxH0ltpIyaRntl
XHw77ulkFWo/NdrRQcNsllWNTZQ0pG5wZ3fAPWaDA0B3gxqmAB8a1btO5cJ4UyU9
b8mba8LVIPN/ABm25BD93dU1oH63ay1gixd8sIIdE1lo45HB8aRZ1QCdts9xT+5E
GOhfMQLRvN4vCcTKiNmkEHslRJ1gtYt/Wgyar4FPQMOe94k3cAKQIu+ew22Rf98A
j6TUDvP8a3upx69yLzA3EEQ9lOgfDc6IqOlslxaz9de+ZGktYXnTde3xNBaLR408
0Jad79pKLVCmJGow4FbPmqG9rrRYJnZta+kOjD2Yi24yjMnoFJi0nqtOx10XFyvv
Eb36K1Mr/evA2M4ToOMpImUIZP24ErpXb43JPoy3Qt1aIuYRdllVO6sgE9lDS6UX
0Jpd7nV9Mv+GYuSq+dsrom3WDE70mUhRVrC3iqStKooQbRDpIK70iGEZisc5qGMO
lBs39XroTSAUAP47CoGdqWwy01OVHuFJeXy/cnhk2UVMCxdjrtH/mM+NEDpULEzA
JfplizRy4Zu7o2cpKAvrooU5oAVtxuNQmuV5r55ADjoSUlj1GcGZrEEFG1Da1aj/
bB4xdEJH1kq1+M1kNARwYqaJ0eP2Mm9124y1y3M3kGUjsAzOX6GnMf2O0eosiAPg
y+6fN5/1mOgMBAXHl5ZJWnAf8MWje+Jt+BFUFVNdyFvialBuy7mRCYx4fcDsZ7GY
+o/WgQDOZg/SgUsxSdkm6gn9QAB9EdhFNNx6QAB27MoLC9s3++ReXUpCW4kgZhHa
nW61mdMF1L8J0IX/429mnjr5ZDEIRVBgS5jqCq7M4pp8gcKq3nsO99dKOJbneHC5
3vbpE4lkiC5kzb4aiPsmQBSn7jq5DYp+ThVH3jL4nwd9mtFnKoJLnPbKOrFDu7sK
HpGOsKvLOlHJwkfgbnUFhnfo0tMjoLSTJhJrf92FAWj8GLuxV/fwwWwABF+yiCfD
XMG0pgAwTThc9lOd1+Ak7Q6dttQIFVaHLMQDvIeZaNYLIx0GewwFcQRXdYkCqfb1
KyEGEO5UtLQC2yHr8qigyr/0YOh3C+OGC5r0a8fQEdAdFrZyCTdoE+u8N3aFwcvs
j1RmPvYPEnbx6/Kt43lx5PEqro818VzvjXLvj2o8cIK1xPCuFxQ01GYhe2r5/W2p
ZwBQK58ValvQcN8YrhBOT6xz6a1bCWEJZzizR44J4oBkr+c6LcdG7jk518WOFmmO
ZmjG8NDpB311Kby5LObvfVhs2eOBOGT5jHS/BYz9bYvXo9OB13VRipUyJeql6H6Y
cjOqRQItxDovXbDLcTVjO6HLNJmr42ybF7pg/Gt9LrgUGLaBX72DfYgag8nDIQDs
8AOD5XvxvktjbHrQWsvDo8f5siR/SawXFO8oqcF1lY+jq+eIZGW+obWTJnQPeag3
bL1cwum2+HMsQAeJS8jYgg5pUpJCS1uYiiWZZTGZGwVCicAtWeCEKQBTAVDyRmue
zGPkdgU/5acACtvYUoIbhmPITDMgSNgKGyInulkwSmOug54+sfQi6LHisjXGofoK
ZldqlM8eMZ+tB+zV8Yja6I87BFn9zfUwKzsNF8oFLn3X+968XaYxN2xFJSxticLm
vBSc01ekJFDIVMKJg2rv/6SC73fuOYIWNBvKTuo5cRgmgb63+VnoQ9SI+hm2v/4z
ixX1d+fd1paTqJ6oJWDQ2JkT0hZRnorJ31tdowQns8iPT70xF09qN4+vx7okARp8
VPzUVl8otYbwWMCEHrfz4pR012kJsRZb0EC7QUPQ3KKQMm3JPkhf1BbPE1fEqt8X
k8shC93aAHfcHPdhZkfUILUW5pRu2UX5hVI7Lkg2dw/o1M/K5PJNtqvIToAicZQB
Yhs9i0bYZSDVqSujzmNYP14Wyb1uuMrK8OHHbWdZP5mLdgkKBcJOfCEaKoTIqKRq
VLVULW0Er9qoLHMkFJR7BCfGIVflwdRKwX7lTgkoaXXZ2PBCwmxrSHFed8NAXq3g
liaEpyb1MFaFnIFEnN9AOApRlQJTvJumx/sJ5RSdcFzKV2/SL/obiEYoQk9wl42H
4wdkKsDaaYsi7OQug5uB7q8Y0TP4ZFZvYU0Dp2dTWdzNVXFUUYO03ZgJ+qhvd0rO
hvfX/R+40+2n+Y7f3ztYjty9qRQu1z6zsL59aCcLiBCaABdqP5e3a8EvSTAQF9hl
ZQyC1TqLZH4DCJtGzoAJIcWi9CgVkFqBfFrGihp91JBv7CQx5Vsop6W8C3f30EkM
UhkaD4Ma926g7gxy4UFKNyv5UbAxUSKc7ZPh2MBn2fy0DNwM9LboQIzckkYNT/vP
WsXhrclYeLkkPVQBe/pAL6dmZ/eEAYnNFBSjsBocNkmwzsxB0R4lVZYK5NHBENUx
JEH2og/aVfZuySOoub0ZYnT1oJSxgKdPIJUrHC3tOTJULDb9uq+45x+FsoxcwpYw
B0sMgb/dC46PkhcdUr6tL7ihubW5F3CRhbI8v6NsBv3z9QwdNP7MpkzrZFXEY6fY
Z8DbwkTNI616AV6Wap/FS9Tk/xbK9O1Hdrzws8UBM5TJoxapovB5vy2G18588Sqd
1xBT4sjbF3bSZZ0UzjnQdJohLLsQiNRQWhkOmvInVFOSnl4TUD6mjYV3lycUeuvO
qW99R96xlu4SDPWbAfgeoJaGePwFkla6Y3C+yCo6Ph/OR7k7gtdefafqVBiftLEC
OiWZkYgHoapCufQo+9S91oUdaSMVQnYRACQGczRogc2nC9YKs6astEYhnUSWPRqG
qVntzE8pGbpt0/Kgg3bT9cvE3Tf9OHib6ZXWOr02QDoBfQ3Gk+J2Fpwvy3NyHP0+
tSHHDmaZ7xe6EXtQARokwAXsBDM4BBIVxYv6NC/wFso3i2wR21FkHn4QrJFD8mxr
elUtxgymqm4TezKT2fA9vFNF7dswUjhp5/ej1ZOj6FuDJ6Klr2+LJ+k9ZjXl5xjP
O2WUyFxw4+ZtOjsecKiYbKvkmDgzkFIakUPDEjkgcKmIkorQOnxQ3LayotOOpsI7
Lgsz32XYRZmEb6Grx3xVN/mb+iQAg3ARM9y418Zru37lP63+Qfoi6GOlnkS5kkBz
j64XNuyMP3my2OfzSaNCWAZ7/Tfa50dYuvHbPYh46Tg28dLUnWNvGnEM7jdU+gP2
FNlX28NzPjvhUrQM56o/3bqR8qKJuqOmusKj76mrn7Cyze6huglBDnfXvayeo/BX
w9ZJ5taFbDQ60lBzhx00NAAtc0vlRAnKrEJy/lSLuMsSR4lYDZe8TNq5uGkjlw2L
GwvNxxC5dDqFBhUPpnKld/DvU2P7jEacBKhaHJY5bpcy6FOfOUCKhoXumOtqiLEZ
EDRti9E9A+2EWqXQPdN+wOfMSuG/MId10CCSQszkq7JxfH8Y+Ch8K5ymoYd6llwh
BO2n939cusAyPzLEvfvVxl8Iw+sprJUuQ2xjiyQJldE419jrWUFd2HVDFGQmtuGB
yZ58g2IWA3vY07WuaIUwrX9k1fP1sf1x4zYmJsQFeY8P8h1Zjwp6pkVh4CVKUt9F
thZsncQyZXQs7QB65Q0yDRq4wpcC6Yx4Cxv3M0f+HcBw6KxKhFU//8u68QUHxDCk
SFGCIiAzxG8b35lnmfxv5C7sTpQxwElloDHdh/JmrCSJDU7rTTAKDFlYtb8lvx/0
+KnKt8rn57lJxJjorWMnQZd8UdvEWRC50SJ6g1M6zsHjYAlB1N/Sm7PEnIjeQvY6
UFUb/5tri8TMlJbd3NjyIHhJ7EHf425TwutA5Maddo8Rk/lPooGbyzn5TaLSQuf9
db7vYh1eII8wBOTG0RMw/16cygiU6WkE8pv/m5FrWpNr9oyqFR0ES6AWZhOZ0Q4D
4+FdJtOBR6XzcWDKM5kcpIEvrFo3SK/hjzIvIBhC9Jl/Cur713ZXE2Kaj/SzaP3T
pHmm+swjupw60IJmz2CeLUwy9pCEVVtzyzDA8hsxo4XKe3n5zy+EeEA/AB2tVOyQ
edXSB7zoelEGZkPfHevVmXJ2JC1KxuOjmXBaXuvlWuORwBG/srLM8y4YlwDCN/gr
ZJLSvWdrbInW6c4LzxZs6zCGsJrxa+1KSzMGVOJay/cQJo8gx2dMYRUxuCsC9ew1
dLQFNZ8Aq/I4taUtS4ZdtmdgyQ2CAIXIyxgoBkV7qJd9vbJG2tIqIwTwk/ZdCAg7
W7xS20GqZJ9ZAgqCNjtpJiWs1lJQDWJbZUQHfEIZoJxRk/xHTuTonR1wSoTRUoxo
ZtxqaT//727vTbiv111bX07PR/ZJ648jQasghhn/s58TdOBXpSClB9ptcco+30G/
S5tcMoH7umhH0FTIYa2N3R+KAn+Et/60iAimMRLLA1HVq0Zj8JEVgnzf9f0CNBHi
yQ10+I5RcBSBKr3oqpq32i110HA9sNMTubH02HblQq9MgQEphsP371WIFBdVWd1a
mgmDUa6Ww5TrxgbLuS4hHUogrp7fftQCG4th0/S+N5W7+enZIoxwn9t5GLuKHq05
Q5Zg86ePhx0Dx/Y6ZbKHoLnSPIGqJPmrdcVx07Q7/Okqq8oQuqgI003jiCpCOV2C
eVSflg1EuwoFVxsvypwFt0NWuTOusyelKkT/Q8FkbmicXLk14n+eRbd1X7zQPJhc
4QOoPoug5fOpeXl8rXgb6G5uZvI3N9uLfjf4qxaRnEGr7gJKkOK6LUIplf2XlRsx
H7CNlPOY9orzNZFGiK6p4QYAzHYQGRhS25/f0fQawphH023AXV2QluDvGtNZkWG1
tRI6kgqMyzUdrNtS/94LCE+Nb6DLLV609VQA4AhwjgJIF0SbmsUnSgHWfKnflT9I
ckFJpZ1FxZMWbg2r+mZ76emfl0Lxh4K3kPd++LLB06YB7KNpQu/THZI3tF4RTuBk
NTv8guyv/QbujUx3FjYTua19Jjb/SnPDpfy3hUEiGaJALEib7Eirp3oBd5vKKybS
3B8NLMT3f1DRhuDSMkkyDJ+li1NRYluUb3illIJwu5U9J146knBwg/Lzp09FYYK1
+zE4BNFEAYo6q0WX52VT+3WrbARa2GcxGDACiEWAoeEde8FBP7bpzQYh/XkXtMIM
JYCGFztz61UCRIkEF+0uQrnFogPUJQookErchTuZVmXwR9YXh52s5iJ+jCyb1jKc
uj88Qe6gxyfqDFjxrijBvnVwycCvrW/orBIdkvKyIPK+nC6x9eY+I22xqkyP1AWu
iesS12TU0irw1f1F8fW4vWyPTkwRbpbtEtKZWlRCT8kHV4QQXptxkOSGL/Pp393N
A3ttsxYFu42SvPCtBxROv1QRb+0QvO2ZAiNLn5Hc6a8gjLtJSgaVU59C0EfLj5Pj
C5uBidkIoY/1ZnSJwkzK1yOHgb3KB+dAXzrTWYacAfbaTe4R0/2NB5xcFxC5FD/X
OpS+BuBpJaB8l7jFcO0DHIx+UlvLokWX9F1OWDHyS8g8rf9HmJ277pKxz6HJdj88
i1EMtunnglA3zsfJlOz66viAhzOt15ghHt4FZuMDOMT9re76AL3Jd7Pn5RdKPStG
ucIDuhuO3NqI+r/YTYcMC6ZYAGGdCzTiMRxHXcq79334SjaxxZA67OUmneyPzDFV
VDBli9eiOUrq54CfEGCmCgzGAUz4BUWpgh/uR+1Uaq/BCdNBDYlCGfOin3Q4LV2N
xByOcx44oKp/16W7gKRWQLN1tLvzn6f935DAEJazzYhaEYUINt8Ddn512YvF8UDO
EDt+8CLW03bYYdQmYdiLh5tVSevYClfn4I8rbl25RhvYATHpT3trARi/4N41eRUs
JwxVvsyn/b84UoJL8seV0Pjqxxi3sPXsXTwapNrVkq3ADp21PJKqmJeAUb1roIXu
ulvTkioZFZOrDweusmRNU+SP6J7A3MZ/BHJWulmBUGryrFKES4bU1ipYDUhUsbDm
3hyuCbQunj3t+A7M0aefzYb6HC5vKLdmIYCJF9xVLBW8YlwIads/VC8L6Hh8mykj
uu5/84IfZ0r1w490cwYYbmwcwfMWmR++otoNYiVy7ZhW0ir2cBzE41MJyXsP/UCz
haQejiYW7G+uZ8G/gw5UYdM1mSIYIGr4XqcEWqIjxKoGkQj20b3Ra3d+CKeANxbx
J6UFlg19+HAmMsKsCi060VUVNLydrJnU4xloqCf9RRNwNm4lt4E6g9oGFkf35Y27
YdSR7MPtRzphwVdn0fEYMv7pvlm34lN09HAmTvPpvshW2eNKPBqlO/kKp2Bt/EtL
0OHvx/bjrkhWM4wzkIFM8Mndz9mle1aosdgO8Tr/vwOhq8AP3HFddj4oVkJrzJOt
jqvKfbPeVExM1xrNG5LTHHpnO9vNTdft8oPNYpVMaK7vTHALY/ELZoC1k9u8IF6W
BgQHLZqgaujK97USN5wFuzNpwKsnpvdAbSzAYKi6R6B+I7MuTRfy2wJapQUi7sTI
gjopl2hZj7r+FE4J+4KmIw2SninbWuauCIZcjEGUWAE+qVRQCvDI99o+6exQENIB
LQ4KVNDejg47nfSDbD5m+EVOPAXswpzXz2coeiHxQg+U4hCCHKNlnzIgdYnxEO47
MEcPyhnV3vUtLrAccBsa292C5Tc+TH2VLwhbo3Sc/3auAp4a4n0Jo+pcVleJn07m
X6R0175AqrLy8NdFAp18dMsDoTwFJXqdl3oqypWgisynM3kIgGzGAzVvIU6ZqIkj
AwxllWTiBJOfP7/p8ix7DqXC4sZQ6ts0jXhbe6asKtoHUFuYsCpwIfwrPxxBHtP6
PHpT4IwJ/UYrn6NRailj9tXxoTIkfHWzfl0zbJkpqXnl6FseqGrd/7NFoJxSLobp
CAGFDixn2op8bWkflLKDLkZPp1QbCX6ndACFybW7c2ZwzaNTkL+MTGgdmHverABA
lBlvsRgojl4We4XlwGu3wanQcpQ8Oi3MyFHwqjvjQKmkUh6XNjNK0xecxtr501yC
i/CEfECNHzudMmC1hjvgQHoVB6wapmhzZhZSykWKSNypzbxBfuM5UE7SIN4feZw3
0TOzfTCw3kyQLfRFxzZLGrfOaGWXFGQlrNjhHN49NKNTRoAL38yF9Lbzr3YglNUl
6GoLjqdXv/dvEJ66eHLroQEp88dWzAyR+mqqhQMENBIs5c72t9CM4+CA7XFJO2Mv
G8GlhCaMxAr3p+vCrMBFhmIoyHtB4TM17a+38bIIVpLsSImJYMd5C1RYGsnY62fB
F59f6DedCmXmCf8+x3TODrv1LICZvVfv7Vk6xlwlHm83shEW+2CytRleC2e7HTZr
ig1sSBZj7/ODTBbqbIvS76UPIRZPVPlixZVegyjQwX152XEsa9P4kn9kjlREGoBP
CWy4VKc2oNeWjyGOMMkRCJNaC5hqgacoxTwaFUGxAsDWiBZbiiGN+BvJidAgrVZB
sOZu/LFCgOdCoTwLI/ncfC7oTEYIjMnDqreOLB+3P3tnFYWA9tVkeTwcVEsa3mfs
MMfYr/eATGus8gjYAL/pE0tRoeHdOyFv/8tq50Ro0Myw6gsPU4vOoxqUJvpZ6WTS
NINsSa8qpWgDPn+2d5nnDWC+otsvPNdnlwf44LM6yejf8i4z/5pwT40bE6jC4rMq
QF6d5zqyXyizvxHfi90Ni740hSe8D8J9282jtWNwHrjCr5/cDn1myNj0ko5iiX6l
ScstYx7uCiFyle6FpIwpoP81PoV2c3CJmJhNos7F1sX55V+9V3kYgdLzaQ/UpGu7
1rBUIIJ8FLK7DL7xWpfu1mjseParTDJwGZ/5QfAHYGYDeMhkQya7aEpKxMplvbTO
mJ4QHenPRIILtTSPxaTqKW5JiOmZglV2xo7QjOUiO1fXsNK6TJeE2ODUR5x4E4Ow
wBW2XH9HjVFExaXMFa/9LMp0bz8KlfRLuvdtWytaXeyXIhTBTouCL6tl5exz9MgU
Pj5v5l0eJ8i/DdnySNPzleu2gEurikMIUOpJemNVD8UxtDUPjKJrOYFdZyEG5vA5
fXfFt6MeB7doPwWr22jW9n86ZMXS0Ez26ohQ4vsi8HXvzBVgq9LpaO55eY4mfqLY
Jo3yS3+TLyeDhXccvtGTu4sC5b1+Y0NlyyaKUzK4VG2kxTpg6lOwCG+Ke5ZUOqO+
T6VIgB5UpR/qlaaBPcwiwmwwlprc9GjTZ+RyiabGTn5Eh2NJZatXLhzhzeLHaIXK
aEJkgSRST6DkQf9FgRNLa3+EhqTkbzFRdD2ylRGDAngSAiDP8MXNzMFx3RsOBAFS
OK989pXml3cSluri+0VwZFwke7l4g42GSX9QiqtyqllI4MKmL27BQSToxxC6fwPp
45qEnjx9g/8RF23JS+4JSTmj6Vmh5N4Wob4DXZi7w7+KvF3LIZ+CUQSMdipuILoH
zOPAwIoXvWCvq3/kS/UGk2UCnxud+/WVjA+dqJ34vO0X7bg6TT7KRnGLMLFHDrBz
TXpM27sl6wEktn7oCOQNS/JQkgmMuLm0Dd5O9t/bqXWQJhl+WKETKZuUnGkblJs0
wJaNITxjJk9fMfmRy7DBMCu9APkzgYjbg0wfzdSUacOrgnoo5zUgf66yjPnYBnXc
oiDxFuy+RREo89x3DzfZppB/MPjp7IJdg9B/WmRZ/Vrb3qgQ2nkCCXq6XEfi6eyQ
ydxu9CZLU4GolRR3uFtdu+ZerrGVJ12HdQR7Z1B21tVrh03hhgSSBxwaHId1C9Qg
Kp8nxpkZ3RovkERVDWT7OFEyKVL1Q/rUBsvbDDmk65oUB5CsKtFC+AQoBCkl+bGI
D5P2/WqkLOHQbk8Tg2qhRSTtQbiNPLLvpz06REcB4LbI2/wadpWL+9v8SKhAppIc
bcif3B6a+gADMdqKgW5YQ6RWAUtRcjglIOYeRHu0OUPAYZHGMakbOl/qq1fBKful
CdTRPI/bPb7mRxMn8b7PiTXeaEioB14pmtKk165tSwZTvi+W8Jv1gRimwKzn+q/t
0SYc3k2ab+H/7YOJD3bStXNLWTUE71hR+1iNTLtSpj6hvaMXUbMsaNJnqgBYpOXy
WTJObNe8XDd7c3xkwYikpatNA71qm4s4Qlr1EXpolliel4h/h6AmLuSql/X4ge/b
Mpg7Fn/3BD0a5OqUXy/2NRjAkU6YupuJOdk5u9gH9BxTIVUQDef1Zo5CBAGZ9xpC
A/D1GgI+BNPQ8YqRbgXf5UJJXKLehl+GAUzggpJTpLjlXYr5zzzpU+7DfCwXNfOt
5TxV+BcZHhsbtylRCUNe6WYOKV7obRYLSvw83P33Tf/a1ChxnvHZuhlng2jBnrEk
lpN3hnHlaHq9432kMenlyjZJyQXObrhSGQNW+8kAf0W1mO8pl04pBQHdY9Rs1nWQ
8gy1huhk9eCe3Xo29HU/Z8euJ4e1PKR+pyoiqspR+N7u+C1TKngYdtvdJkG8Fv17
YTpCbTmXkhpAiJGEXvvUyoRYVHNDrOYYq1t8baMf/bqrEa/RcxZH4FsQimweyvaP
R4S+nZIaUXSiHrVlKTyeoSzp7OiqeU//yLewdkj0xdjqrQE3kP7WkffizpnjL0M7
bEDy32BilP3tZ/H65J28LQiDxrFJ+aXjA5QXNbN4yyfjwAXj4YvizmY2hwhm6Edj
lSqjiagooQm7WHv5uPHc3GEQWQUWLn+B3yRQn/hPmNJHF8bZ7GDDsKukvDdBsssi
BJNqEqJl1IiukLeisrB0srpn5Wp4KRzmL8Y6L/KuMaOUgPAdZ3hbI0cJEsGBC2hK
kDpp76yR2ns4tTNbPDJCB/MsIy1PvayFeq65fauYmhy5U3Lp314KcMV7CpcqizXF
xm/pYIGQ9XtKkjqGi7+SE8nB2ouae4muknr30UtQwpi9ciALjBw4RHrn9GXsjcSJ
tIIUrCQlJ/XPCiQvyfyoaRW0sxz7zF/HjAV0m+2VyPSTGu/BgnYUPw2YBmhD3m4O
7/vyP38i5ArPDw5yCDTBsPQN5si/UiTOZ70G5bn4FJg0pKEEqAFkNmcU/zc1IkMJ
GDVufRMG9PoKSQpEgyL/k42hPx4jPhi9BzrYuXKkonwD5m9FUyYAKy5g3xXi9fA2
iAXizFfupO3IO6ER0tMPpdJToqwvZSJSRgJO6md9lC5etQycTaPJZdHoQayW/hcu
JLEL5P9UObsdZsB+/eb5DwERHQ05kpxvBup0UXv8FOgSYDuvvGNlL5Xh1tDiUhna
mB6D5rl9QVgKUunOHjOCaQTMz+Px/H01sfl0oV7LLTrGfrt8lud7ffaWJHtCFKgM
ZETstc9rQ+KQtQ+eWhB8QtcWgcYTMjU69kXG2smytafy4bbKvmuXTFCU3bzbmSma
7ytS1xmhO5hS/rDkkVxbr2yp6tWpTek3SowEf6ZVHMKp3wdxWrZ0Fxvo+B3twMPY
XyI8vUHpUBHIWB/PAmc2wncjev0LIzHga8q5hqkEy19ij1KJyLMH9kMaOJttu+SY
KJSFFYV+5ZC4Ll73q0u5N8gAueaNL1JgtP9MF7us9Zj7/942Wo1m2ocZrtUwdFZm
ZpOcaN/j04c6lcHvOrvwBtNiOwAI1YUvlR8jcG512dpVAeRQPev9ahQBZDsQ6xER
Ljmk8OQK3fLYDpTtS8sqbo1k2k1W7ZVjPiaikXwfHZCNHK1hRowCDcVLyxH1L5Ls
Nv/R7LQsSI1PoxI6deF1LGDr852mJJAoT5JCssF+P4rjF95FnnUe7BC17rcIMBs3
05mVVzb241DA7XtPszGbd4QxD0daLz6uLHuWGdWmTFPC6RL+kz5c9GlA8dUh32Ex
PY5uQhhuhqqftGomMS+gVj7hpQwOU6ANpbI0/68VQPLmvTtpUP9KLaLFw0xE8Lqu
Z5APB3BLFxycz0WhPtmXdxvtHwcJF2Z9ruN8APg37WKdtvU96kVekfXFLagQDZoT
us0wo6tizRk/hB+XyL2qWDEvAnQUI5sPigLXIgZIl9TTu5FiS0+GQfy6s8rn61ry
0IlimuR6yFpwqY3ytrnwQc4BIWHKc/XyunL+rljNtGhSeN39NjDM+4zM8P/PdE4R
Fq+GMVjW/Tshi2npRn8SI/7Vutu//y+kLAtYlceJiwFxfRR6ZnLqcsnpsqlCU52h
OWPxjLBgfiJE+19LsWD/Hgrcos0wq39Q+t7fokuKHjYyiLwS9jUkwGHpc1mRiNiW
BnSCTCMFckWefq8r9XLufw1S+35p4mmNBuVF4tOoIvP6lUk1DdGcrQJXSnynFCu9
HtgzVPktmtBTqg4feRkjH9brk1G2gGC2VvcwXg0RArbNj9uVZtWZmo9zOpyV5sWQ
CHuj95h3R4+lhQbNBPqt+vA/0n2aCK//u+XUbdDTBEacXgdm6OuTBi+ObVB9FyTo
5Hab3sX6/5KHbuYzZ88Zo+d8cYY7dmhWCcZVyAuY8ILgl8oGhMGVCw9UKTqxIid3
njpVCXWqikNj6U71FdNhwkaVVjyad2QvPnsWHPceacSJ9c3QPD8f/+8jbLEm10dg
VKvmNM7ysVbmcWnt34EwCLLMx9R542yDAEB5HbmE+9tZnibXE++BfI/2M4/bOHBw
HvmVlEuTdrtamH1pG9F+4ioz4NlkXcGV80/q7cUQlwmhUNBmgcD1ZlLn7kQDTj4z
toEEmVZ8S0ra1X27emyUpHjbi5bWnxy0FYS4DOqOfjjRmRsfpILJS+TFJk5tPL9m
KlJmnW/LEIlapr7lako1YGGTDemd0xHK/0AAwHIv6qyYW9svWzPVI4XTqmsNPIIq
c5K8mzY7mnBCCisDxmnZXrZv2Nlq2lwbDvckYP42OzE0Iv/sG770AMgo2Gfw6liq
ToIp3IjR+XDgBN31t21XQaAbDkVU6MUVBnIVwV1h7tBV5QFTXaAKvGxAck2NXerh
hTkqoyQng9c4qtZSAj3Dt5J+9tz7kR4K43VT//wbB9UELITfBU0nWohyP7aEOAnK
Z2cyr6MqjChfotPuniJBm+uyXOacn+flsIT7N/9TdabJjdn/r0cefbC1pl4la3d+
iElFGWXXeSo/2jEGvJC94QT+3nWDaOztqcgRYASv4zQfuoxVAWrH6xgoQmINklCR
xWr/FoXGKSMznOe0uxxFo45s9+1G4cBGmFDoWk9ndHC9QVRSUMyDfTPF1fJGE6cK
0aU0fRkyh7LLwZgXudLDJXXNbGovlrnJbmGVn4aE59El5oyd7lAuOhHTebtq3V+k
AWk5RPSamP8qjpWgV97W+wM/lac2EzVsrpeXRYBTPSK/AdRgu9/S2MI6IOfeoLmm
Y3Y6rtUwwLCF+u8ymmJb+RMkgryaTjA/NVonMNBDJlE+ObDvVfgBsx9V+Xl/ETwN
J6vRwqzGzuwfh9CnhIR758kjLL9xZ7asZFZ7P3vRzQSks1POYCR0HXLdpfpaiUkL
VRqduapvl9o7in4tjdI0MRFOLUI90tY2TW2GKKLHop1wInWUBx+K8SQioAzvb6s9
rekL/v0xBc7cgGv+EDldntQptOc2Up/RJnTfe3nEgaTzIggu3pSLi8tdUIRH3Ld6
bB/BFKt+LoEdmQPzI5IwCWR/K5opV6Nxoq8nSuYa4Je01/E5mEiKS+ZFPXSpfS4s
EYKkUHJUbm5b0Xn1Z2whFgBOvZ122X0D0SkxJArax/sxiou/IQpaZaYoird7Ou7F
h/LaibWMI2VMkObXyErBcqpX9/yqw00fmfzTiR1A7zMGJ7GIQQ/ocMKZI4G5a+sQ
/LufOElPgEtywe9NulK+64dk083pQcdDo1Wn4TFjv3fPP3ryn9WimkRkrd8pR/XT
92FxjzmejTiSoFtEVsZV73YlQxtst9HgWK2H2+ODqXiqJnICtJBSNJpLbph8Zpaz
BWqRHPjNYJv8tZfzHygJ78Kdlmd3Egn+BcYoqH0LzNGyv339XhosdiCcawo8EUQ4
MKBG613zVeVcRfLrgjn2jam3El4ISwpJWg8wEG40m9bJ/fSg6JrEk+TIPnGkNOC4
PetNb6pGM8ckWLEhexoIZ7sjUYOH0CRowymPqNUZur5f7LBede1v3ulBq4sV9R9W
X1pU6GfMNxk69ApOplaZHAhel1k4jTep/2xlE/aq58qOf79gpeyU5btNQ3z8Thzu
WkzhqZgBU/89jgWbvjU7SNed2COKI7j3U/T4+9Hav8VuIvCk3nbrxS2Kn7/DpGeR
MQUsdfRhqob17mxS8fIqOSa+SWr4k/jsBCeUZwvJifyuANxbvRfQyssSIqznswxr
CCocoR/d8BIBwaAlTbYz0wRymGMBj5MQgjXLFlVNaVVeMSK6RxG4W+mngxvfWSji
5RN6XoiUU4vMszwT9KYu5YTdcJrA9KI5Ihy+rtOcsMXQNPw3f/HhkRzVj3tlT8TB
1JvASio/fklKPLkqlEQt9OCfFGvhZOOUoF39BxXLgsFgXEZjIHkf44H84/E6P+mV
DcY85Nio5LIQwg8qGmbetc5jpmG2CBmamlWUaXoP5rzBs6ukL2xrpmjLF7KMftOe
vnteumgzNeUJn0r/G5yl3J0swbmZIX+G61SrWbHQZTHKkmhDL39RqFEf1jzDV+L8
13t9SKfgrbtxi+aEMdvTAYFPZY2PTMb4CT4ibXighDzVE82sS4ZdEoR9Ry9vz17x
8EOrdV8Avu1kPPCAVtZLeW1Php/rcyKGyr2RiNk0qVwp0bCkPZ4b8NxRI0w+vjIg
j4tv6UnJaong2SqrajVlKeU1O8t0EF16ehTn7WBWoXXR2wTPwfDohFRwL9m13Vo/
85OavrLjPuDdHx+r7oTRQTlBPPPgMFQ1ElhFx8lkA/4e/L7m0RIXuUO9p0XeRNnH
MgSCH9Lc9Q7TVq6xP0zkgCf0xfM62Jbbul0QK2G3imM3k79vqmN3gDZ5buQoVM7N
lOLwzyWRzXsKUF4dC0+l3qTR/eJiGP3HG9KtTEql91HtRAHBE6lPj0SsOAUZ1JNb
f318O+qwrEitwQRBzU6CnQgHw6Lp6CYIfFb+SnWdXamRofsN+RcYP82xeeDekp14
mewsDK6e4PFoLy6Mp5w6v7GfP2pMvOrtnszpuEyZkgCVWvPM6yzgIAUwiyLiOS6/
x8m+qxOR1ytPLC+Mpv8//slwKkhaGkbdITUQ8xgWR4V/EpjOWYuPI7zXRkm8fNM/
mCvlFMKGW3y9BU0dlyF58O6F1dEDFfMwaHlaRX1VbnWV0mdkVsfYNTy18OcAAxL8
ZVOd1+lglE/FcC3Fxl4X8BIhR4C7KodO7hwfVSYfsOU7C+fXs4K6PcFS74rUzF3m
GVFpUk/pY2pxX+b+fMflLmZcX7sp0Bx2rsyWrvYpAmZz+SrnWaTMdAaJkXrZ+LPV
t5W45GUIgC043wiMKizepbbiHdLJzyD5iFmU9jmen5mSpQn2vPhKXoLjdQ0MTnjb
mONFmsZfsL1VDSJCio+Q4rE4rSXY1W7yhtDbP007AEVSFAdf8M2l+LdrRcKrajuU
EGF/cBRLLcxhx+UZZjrT7q31ezpFh+ey+M0rJC07AStZI8/2yvtUkvj+Va52pG3w
Krejk5n17kOOUufQE4xaCmJQPtfZwaSJUxKMsSxw0p5mbSpOAzTcO/eG4YN0lMmx
uU/8lleQ9MkpKnvudeLmxF3NRktCEPC9M/1YtwGfo21sYFgx+qgkNCkfCuCPLabT
MQOPN0JGIWyqPQeSxA2UXni3iMGzjiSzBteWrv5KD6VsG0Zo+6NTD3PREE0dU39H
5QRpjDT1ABRN7TzTzTEf3hcOpGRY6RA1u5WxW835tBLpBB/TYgOzcxA9X9yfuYeD
Jyo3G3CB6ZsQdAGcCNwZSGJFQMDZOoRWrzVqUaquRREMUBwQ5ouwuWoSODYR1swy
4UG+2n8enCQsdcBwIKNyttHOWjo0nHz1rx4jAtCOgThr0qzyc2j/BZ4tzFexUASX
2rtNpol1s3jNocn+YGTTUEvP9m/YSkXTlSqJ7YMERMTrl8aH00/bwgVhWhkUYpl6
i4Kt5pmWEeMjCxF19DUNEkL/mKgd56s5pON68S1q+YzE2qHC1tsuLaqH6VZqF9W0
gFhbHT4zQ7/UEm+/NHM2P4pzbwGhe89smI7eIRy0lH1J0SmIc7Lc8qKkm+D8K7H/
ghnkIHqwBAF2muVSmLSmblEsY9ksmc6HeGtaNC2tBLL7/E+icxjO7AVF2ySupMbQ
ODvCsDrJqKPWRcs2Cbqwh7GZOEuQbMhl+a6Bfc79CBfcNIttRgfqo8bK4h4CDddU
0SwYBQH+xPdWfBuWCP1/SgZqQJ6MMCqlrotuk3ZHmSr2hOpbLOXK7jSXMzjpQUj0
6tX5QGv+ye/ZNsBDHpoMxGM7hqEY/Tq1HKUH4LwrBIx2N4hcgi5y1IquAk8lW+MH
9MOqeaRtWY+fLf94nC/djNNYR+efnFMaGCxZn08dV5vKDXaEfjncnvIiQ2hi2Q2y
Zhu7Ro3VJghtCY0n5X5zbuFVJ7y0f3k7cnILjIbWGMUZ65SwBtrCbLzo4ixcTDJg
cXh5AiidU3OqrSeCSmXgyzFpapYsORieqHnO1zzOEYP3DGO8K9p4DR55lH0v62zo
DED5S424touQieWRcGy2EVuoIjDBDc4kvmQCBvdH0grPAp0qnwQOwa4PxnbX3n9a
UD40VQzOHxHjyw9AypLz4wK99EmcWUiBBKWchW/NT0SSDiP9wgQUXLzTdtI4l94/
3eyJA562eBRnmaDQeVrGZtYtnRlVEZIZxJYtGLg+jVaqdXU0MLHlBeNeya7hvn+W
mVsqrBVJN4VPJtxJvY8amY7uU1sEVQAYIL1WJq/wzDT5IMkxfhWkuoL3nc+kr3uR
1t3wWRqWNtoWU9p3Ug/QugXUEjjvcdzF2pu0+3tEhOIH2RS7zZvDHh3kf5Nz8ZDr
xPqVPzO+i0ySr1Hgjw84ev3SyILJ0zbj77GDe/u7REqwbBjaiVolUTIwwkkiJATR
43GC5/yc8Tmzf2QcdbHQcutamJ4ufNsWPn9m4KBhbO/YUnOSkl7LMLXRND15D7OY
jL1Q+z4sThxz4mJ24F12NYzIZW1pACyCdjmVF0m7vq9xF838leNPp+Oa7wo1Mr1o
vmIAdEpfa+cmegqb5EQJaZ9ImkmR6PSILa7w4WfD5p/EgFlHK+2r6SdGOcGWr0TE
eyB84hMoKE5+Ma7mVBL1+zHuZykJp8NQA1qhrfyYucE260i+vIGX2KZfiZOoOjnb
wd5I7OjAJdt6AMdmDW1x9ZRRMpq1Rbg0YYz5yh6Fe4WyuqfnhO+4C8dGmEVnV0t+
e0rxw9kvGq94B+JRYw30fR04emyuxGvYL3Gqi4WI6IsCVgeC1WF/an8Or3vpvYKO
V7e9xb2T9K+79qXl27URcOYcr+FWpY1u9PvOu1HtvVTMb2+bN/Fg2W3fu73HfcQ5
5JUtzu38mu4FOJ2P5I0hK69IJyj4+RRX+iAWohw+U0S1yYdip3yrTAUwqxtpsBFO
l1WvE5A+FdzVaV9TqGKXEkKbQDf9GjwfbYtmPiC+w9mtYmAP095/BmE9CwFi3VVJ
PkQ9REJCHGeEjbDMIOZNMYO2oZMG2BZ+RefKimv9wbmfFXS9TjWIrOOUO26SBPet
iRcw4SXzv+P08s2vDYGLVq8sF0Og+XvNLK2+7rMifQJbKQHKASdfujOSN7uT1xmD
C0HzR42NIWKia1UZe9uHmD22nGUMOmkXX2m759NQh+CDjaiwYTuNArsikU8v7aCA
QRqBT+Zh3ioUgTKutid7pV0f6Qg7oFynFWaozbzbB+GG513WeOCY1XhH8o8JGGPa
BU32kRBYlNhvhjz0/wiTBlAHeB34/HDEsQtHizkLc2f3QPMaD16s1zXbR3QT+uEw
+FjByrIbIwB+zivI4dWKe6NysBiF+ACLicE1/yZpPBHMo9NsBY6zMtiPaF3rUF+5
VZHUz++kiurV/oi45iIAkoHbqaSJE3UE9eCLplvPygYWKOpgAmio003mBetd+VuW
ChxXWNhLYEX6pmla2st43hpTtItTxpMNos3nS+DwvIqNs0hejneijKzjesSqCBbR
Y1KibcfKrQxFN4qGR0SMINKtcHZfWUrmYLp539oQKWOy/iqvkiEJos0gbKTngC2Q
qOiWSZ5RBdCSDDoKB0rRQkM1p9M3wWA2dkMiZsaXNEs2goiPDw0RbGGfAkrPABI3
FbPW8gjZARbg3o/qUMFoFFZjs4ijfd0UNXtEAuVL4SNWWIWrK11nJcVHWIzY++9c
M9f3HcypWRPpRy9K8R2qd+TReYOIgndQ2zKa4Jd1ePAylCLj8IDdj1qqTvb+Fge/
gZuETFkIuXj2trikjrXe4LwI/+9TRVGC4zWr6fChOLAkXRJrl0752nI22oYXTAHC
PwDH74aJeLkfdZ7bJst1MaQuFGZXzBuJ8jxjIQVGMzJ2oIxiEIYwilOC+6X8H6v/
zLadB2JlgUOAY03pyMhpqF8lSYXmXRVJOHeN4/gvGMTkBoHSBxyK1NlfZol79wJt
5XR5hcocAvaFX0GC0RIMTnVV9RnaZtwd2CPLPEmXavzQEFtB+BB5siaxaYhp+CvC
yn1cq+a2XHx2XpqzWmgMiE/ygwdHGm5Wyyh1URqPQ2OpaW8DdIXBF4XwGg4q3Nb2
BKMoJbmL/QopVPFMUXFhYIjJ0LD8TwsDefFsx5MkY+MNw3wDPkmn+3m8BrYbk+O+
o53R2mBHPU6NnQKgFp7mm6EUmLlgwz2s9v25ETfUpSxuT5QNBBrcCDnER64xxad7
3CjGoaHwoQNQHnBAOc2s/An4LjB1qELa7mVmhRjpPOAk2AIBL4IueTEd/JxL+70R
fE2RKsyab/N0Hj3MVJ4CprrfVSuTA6Z4AITOw3H3MlJWRxvMnIRMIYaVFCcyppiL
NbM0dQsje0+k3Ny1WTmgqXEjAFREDQxS8Rwee/NLmykAUi/YmiChxY2mlYnKuUxY
6IKjpJRveKqDGPY0LLdoJqfEH3u+bDiyqD2sQjduVmRGscWVm3QCbtbNRwIqQPCc
caBMhMUL4fuzTCtc/nQBjxhqN15karMLM2NDySb3aPp3nt/YavfP2IYiBbuVUIIm
UzDFQBfkxBhF7pIL2sbLW/EgYNp6c/YLgOzR02uh7kXE+PjeplSTkJazg9uISNzu
Xek9BSXc4+7p6XxLu5q7if841Jnp+B2gnBwGbznZyDVV6bb4Xh4vUe/aFh1MgBKb
Aom31SIrxlcllgLEYUok8/HLnyWfiJvRhcOH6Mf+IJAga98XR+5SQlVogP6XxLsG
s4ZLH36cO/gcAk2tL9fK74xWCPhHrf73+MLjKcEaz94Wkqg69CevStcoGRvLBmRx
TdRLh4v3pX2UIrOkNPfyyuROffa/VRKTO/uvxGePND6TJDL132IVQVEesBvHHQAt
zOxPf3UildqEkE31pwl+krsAFD2tOHH7yiXUb6XhtWku2gjtA2F9+YIesC8Rd5Dg
6jiHE+YkRLDAADVRbVycWy2BoVRhKovu/h0tn/mFXUbGbDlZjiwMumFMhWDg5F3f
z5/HWR4gCea79p8gzwMBWO6JlKkxBAJnKfKPzpgyhUhZurMMKkMAVjBPpWjMHI3A
2n3pZ2U2R01rIvVkBI/Rwm5QjjKfYq4aMDlKUUEyH1WLsZgMrxrTkT99tTMqmEYP
gacOnH3kuWwC2Cv5fx/pXnhaQqJXbAKQrRYfHPV8QPUnt6yDT/Gv6PN+6yyPE7PT
EiXo+/W2bTrd8VtAUxSu5522UWm3zFsKE3soRPGx1WpntuND+SBWLEjN9ZwcUKQ5
dnOZo3XGZbNd0s/KXW/5tSG52QIKBptz37u0RMJ7eIPN4gmMMv+9+7l8ZFYZSeft
XTyeTBHEscVEM1CSzxMeBS43vuSQgPts8p0fiM2A/F0=
//pragma protect end_data_block
//pragma protect digest_block
c++At6bp6hfzbw+LNrTDElxU1gU=
//pragma protect end_digest_block
//pragma protect end_protected
