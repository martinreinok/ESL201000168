// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 03:52:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tfLZ1KmhLZoNhTUpkRLPgrZinyij+ZISUTCrqDFFyM/3ai+3m3xxWOcbH1VtbuO9
KVlfCnbcpVW9Dlb39LCLMbyBLS0gUQXWkTluiQHoLgMEnJ3k1k20QC16zbCq7eAm
K4IJnSqUaqHTQT7S8vW8E6BzQBNbHnJXXIulStOmFlc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 38464)
W5pZ41Whrrfl2dfZI7WD4IayooAsmd9PHLM+wBdSW7URyvIGy6f8vvODvPIZmzQE
ugIyNvYqPTNRG3yiJORvoGvLZmXpX/RhKCcbFHOqYguehDmVNFFIGSqs2J+SYVHc
uhmy4VGCGq2s3qq9tWqtP2fKsUHiznRTv7h5eRYxV6Fe3GRJDncl1yGzZS88P5vK
X6r6ZBOUwzRW4YEYw5IEakCRBQeO6AhWlwqQ2kd6dbauDGzOVmzZIXPr7PxmtIgP
8AB1ildDc/lCry0JelsocEgBios2xMHuzyQEEUp83giyyb1wNRwt8vqhuzfC4eRT
tQ0G3SeeFKUIU+YcrBkpramjo0PoO2xUR/ZPTdYGdwRLP28RWl2neUWGfDvfKfHh
cDivKwtSk3/dVyW/JVOOp+R95+v1VzvangfwfGeBCJqV2VdUpioL9wTZQ2fXJ/nb
z5vI1z2FqvnqiykgFDr4+AuKGhoxxVdiutlUo9qzL0rxypTGJ7UZc5rTC+Bm5sU5
RupQ0z5FIzFuQe/g63HGObhK6EyTrYqwZwJpUUP1dOEXij7zPyXW6uewWflNacb5
z5E6GE5dOYTRYFCaamlXOKbk1p4zpZjrLzV1f+ry17aDYLAYubHDhFjrFD4wJUMv
EqUi527FLKdh3Y94dR2vXST7pYsGUyhmT/R/XQipSuAgy+6kkyr0XE3A9bFwBYue
NhBY12QEz6mT6qs5uTaA87i+UQ48YbUS6UJdhUOqNv5nT0uI18cr1hT7E6CSAvQM
pkqqM84cD0egcNoRFGMxB5L8R+WRbz+FPjHDMMgkXDN+c2UWPxp62ur+lXo3XCFE
88qzfiYvhxc/58fPCA/Uy5neKmkw/gzQNmUU4ia+5qRX//X90u9gxm9QUNC/i20I
idZt7pD1lLJur0+XNJEB9R2TyJ1TMhGhU6ReRMGNeRW2XeYEDFZ3rwPLfAoc0mBo
dXJNJjQEWxCRqB5fkeUg0c0LnEDUtVnn7pdDnOOficn6RiHUTSt+i4TdTix18vkg
RPCHu53hbV27v7KwvgBxRl2gIEB2QpacOqsihOeTbmmG9Vw+YSurTSVlLVCY79CT
WbUPy0fsJFsTbJoBQKFr4cjl3b3iZfeXKL49KI2jO9lVH5l+o/KPBaPCSmQ9dSwk
BnO8lFT++Pwl+Bmh3WeDGB/cO60mwik9UwG3WPnaAsJf2FfGnMGFDDpDopt3kZ76
+sEwqHeu/5ppCKBQ0wWilljJxwI6gBKCSauf0LoaaKwp4Zaa+xKcOLSw/g/rYgho
9mdXAXde4dFAHvmHqB0b5lQrIjoB2p0sOIEN6KPYkgVQ6wfTfa8yxulwlXNYfKqg
h9y1BV2TL55p7oXUtDAG3VJzx/wCCa1ghhBovlUPPJOZpRDQ3son+YKmV5O94mQq
gYwa20COVNBXw3NIgmobTU7j8KSe9+SVXbx2zYVKXZ4lifuegiG0t0751sp5/uqD
DjWbsNX7cTXYKo0Dm46rF4dnd8s+8CUQoC3CitEZx2Xd17MS4ULIU6f9/kyWWO33
bOUFgI+WoSykj0kGM9sa0LRRbv8v494whTEHGgNuDR5h0BBRPV6/+c90MzcSlahw
G08y5KOMurGA5JImBQhC49aGlTF3LE/MJ1QK9uTt7H8KOkMBT7GDPtsDZkZC9S8W
iTxs7D2pnup4rQjcgHNqEm0fwq56liS23u79Vjztgk+qCKEcgMxFY/aSmiPVQNPT
iSFTvUwowXdDV+udWO4oK/eVrRvuK3KuTNaVmJNEa6o9Ib7ZsfOgY3Iq+O8wLLpP
0xcSNy8cnaz5Qfip25C8ta/LycSRPu/WlrzmalhOCnAee3qqIu05sV2gzy+ubmDa
NkOlfs1L2121S7mo7eM9a57zqzgQu6teM+vnx2viJwu0A0fSkJ9jlz+BoTHqhaAj
rOA8gbAYDvbTbZq3/rOFy3JcsWEUgFc6jpz2Wk/KdknC+hW+vI2QtyTPsMqnsEbQ
8J0hqeDYq7TIxLujeuH5RWh74kSOfsoCIxiZcghJB8lobeDTO3ZOVNRc1SS690uC
WyboNWXrpyH4v4ErS9kGI/u6OWrhk6cg4/80IV+3uF63dX4pm0P5H+6kh/Gzo4fh
9nT4mDiq89SyXSsOeTf9goQoag162Qz0qe2EHU+gd3aoRrPvVPJFpaMjBFlwjBGz
3cPxxH1tPESaJneGbnHD5rBIduNA3vkohxjwKeZqDJv3aszhT81elgjhEVtUaT73
yvo9PN7pyzQ6kYEO01v33js+4TRPrgTQkSelAz8oD/qDV+kNb6/NYMKqOQsNzIaL
8AlZsWLD5VxpcImDmkNGDfJIIDIg8ojA6WjPx232hu+TWRR11knESdUta4bTS0TR
tM0cvoXrhQJk758CU9QG5v8hTxKGX4NXtyZKW3rTMV8YdTZVUhwpViw9BQcJFMcN
zS7FBFvslHcBIIaRiyOKbfVM95bEEpExkxA/OlwlwcJzV/G24UVrEJyR7NGsrKz7
LGfYVWL6HR/XHDHxETDXzRgGVMDJ9r36q+OUYwcHWybqRVKwUegnVH1K7z7rGDNt
sZNCPKHqHspModo6aqpE8AZmzYVDDUWyI/a8armNLkpUb80No9pkpFSbUhxtLms4
r/o+7Jyz3tnr1tNyf2F4kgQkztdyl2BX2rYiMy9Z31BeaZY28LtDQbb5gk96MmCP
rUReakj5uaIWn+0ve4YQDLBiGZhgOa695PYnfabfI2CW4mNJOcqBhqyQMT7R3/lN
vCqAfxCOYATqXOBks2S6+238uYCfeBXrERaRUq3tyAZ0xjAEpxsoheLRMioKQYsJ
3H8fNeK8ppQ2Vcfab27S575a13oVuEAgAm8FhORMg4RkCehXozttC3PHhvlMAwwW
K+LStP4gQrRay8R584c7SeTNrik98WOnS/f3kozCyQEf1Ja3JwDeIfj+WW19zPFp
9mzvP1rJSnv+Ox6Y7xb3S/6PAbrcI9bDROuBes3+hefn1dRkfVUfMywttFLgAQhr
N9BM3YAmErrCRyi2o2BXLDix2mWQRU/8djdgNvGQRgx2PMyS4SXCXd570llm7PWI
oApvXULxsl0sjN7eqi8wksu+/PX0DvEd0JqzX0adBJOs6k9kAIBffU22m9KN8/qz
72vvc26oA432KI4rwXjdbWZxivTPdL5Att5+/7SDSYPQjpuQNv7q8NFwfxfj3Pwg
SppbZ6/0KW3GGAtor4P2X1YWP1ed9Ap3kO6BkWsFJodD4vmdg0r/Wgse6jDtCerx
IsxCMtvFHJekFpDb7ThrvZz4seDyMoqTGrDMUVD54BsSh2Ux+iu9E801ryB2TSws
Q5Mz6M1CZavzuKPqRFW5RvspPBcfOKmQQ3Z8OlvtvW0CzRhZdpgVCw7kAVdzLsba
nCd+Wku5k+VCsymZRmba+mWLfmWvOlaBVCe8TqOIKQ5wrwHwVzOSdEM3pmVzo2sG
tb0kw2PzAHfSDJan1KMuOtdBKqxiW8MDl488TC1NqGTX7yCENO0yPWwe5nhJO6kf
9Gbaaq/lo9ztUHwHAjs0mPuz/yAz0nCvyH3ZAKR8Jl6wTvQ23iPHfYNBaIn3r+fD
BRztCQs3vAl4jwJsrJzgyrVlHna6GhowrOdtl2KelxrjtxrMBuybIwMp4R7l3gU/
vCb/iJdmxV0dVsvkYF9y3/by8Zl5qG7SUt3kFDH/JzdvIqVdc5x3zE/xp7t/loZw
nbllR6NnxZ1ZhPUNgCtpzSR1F7jexP9SO/uCOYdNGnZFRozEWX1dPQQNGXbvfNPA
yw3MHeT177PkFPcz+VZn2jjIVrK8O8e25vJ9oO844UuKYmWtC5j/5r2nPWJKEPsu
zTDsz9kZgz22WMGhBXdp8pbpCO1YWQGX+2pP4UK6jhgTp5y810KDdTbpweSGAuOM
IFaX5NRHxOdbg3KJiPzAx4s3nn0X0HGLcYfF5LlzRq+b/WWoFctQC/UoOZjdpBGx
6Hj31NSk0qpZqI/vzg2A/jRtx4vsMmA06MzS4HJIzCWO37FY1KrK3eYwcK22zrsh
5+7Ov3XQX/SaYB+k+vIiG0RZ00cZoVj994gyIbYLliJl8Y7jAEhR9LNialsn7jOQ
VIUOlHTMgwWFWBgwZU+SjQcurKHkg/YoMEDK/LHc45TxfbK6zXqhe+1FcjfT1T1c
UpyCp3wHeP2XmJ0zb68cj2cV3rPbsiFALBI/dVhqicwEPE55xPHm/3b5esOgKVXo
RCR++bLHudAOUeADLOZ4/4+BVJXWahbXwRvgeTwYhx+TzwUXx8sTE/LsZ+Dts46d
SLcMeZtlpqE96tlW+Bqqo0HDj6abqhI2D+ASg0sbeNtIpAOfKDPGqprVDaKESXR1
MboKwUd3prXJR9YVzPenPywFP5VJiyBc87wk+tG72+BShPTy7OmVr9CoM4IzeEia
uFtw6saTt1GAPodOaWYeVx291iF5VrOErqU85tou+0xld/b7GcfX5+i8yzSjZEgz
/L7cXu0eobmNaA8cWitbDBAFvTxTzWLpv1CIQ7YfWHvKcsVRXNNs7wLiC2X9DHOK
0TsBsUQCcGZxSYUxZwYJpbrrWLdnyQs1CtWQT7GuQe89oFMRC6K4oybDfTdjj9yi
3n9tMuan1Z9Xc+gj0zJSTfHt/1LtUF+CONd2r/newkLlQxiUOKMr2F+D2fRLwi9T
m0D+ITmZvCHQQKtpKXOKMEURJoxfT8lu5wtBxpGjl8g8Yu2LvZ0nS8OSJCDbVjFy
T4Yi61+0O3dLMK5E2ZwbV873fSJrmoFdtfJOUkFkvNKX3yRW9Q1i8/cHMe+KZE9A
9O2OWty8rUJvtx95JZJBl2FLci0pqUfFNryKzCby6hCq0nEMQpbdesuNDpNRdKzW
7E/SPgpvhlkDlKvsFhtZFYQlFhqaBy/0fmXPbMeVfXr+wFGUO2G6KMqGGqgX+v3U
fy4/iULeqbDokDaVukA2145+Kf9dtwycQgSuElCujI0MpNDtzqhaIH1BmxcFoV8q
jSJBpqZEd7Y6W0kJAOhuI0CBFRrDrqjhz2C9g7uvnLKVtY++wAaEVw1yv8fTbDBt
5s12XcowdafIDUiAEjgJZM/o/IaDfDu/vRVbkj5HiZIh6V3hBW1uS1aG5orzqIvS
gXspMW1QBZtfdqkK5v/jZlGFDWcyv5FDtdSRRlHgcOH+TEZ1UiDfuDmAcEGUNT1J
T77szcPKmOVTmZ8qTiG1uNGWT8b9BlBl4TasZaZY9Yf9jtLnTQjk+872SWDWef4r
bx1Je+B/wR+d7V7M6zav3PZtj03aEnbf3RrT08YPgLvCVXibqjOUMYP+u+Ou3A7L
hCH8BxRNr0ZRN4Iq67HWu7bdq2Xpp8KoR3aSAcfj0ua4nY8/glth8QzOHsRTNmIq
jHW7q6c5jP0EebpPtfxvBxu3kPPHHYx7IbdFrCwpwjH95lwJpXeuRFDS2kw4NNCs
bvdT9abf8TiUtAisB4dK63q2gILT2iIzB1ZjZA9CA2/F/JYM/0jmZMMwyr/cw7cS
EMscy65rKebLAVD6jGoQgtAp+0LJGDigWatLSJ8JtQP3SeUH5vX6SQPjm7irxIvf
UOl30Ka50b4HEAwrDoI4+xGEzQk/16yxFXqndrDN6pYFJaSmIqa/SsNYPeZ7exn/
LP85aQOX/1jCAGuJKcYEeVEAybKvhi/RDQ0JacXCUZ6u3SaJRB0u0CCO/5CcsL0Q
MF6TAvYMgktGa+wraV9o2aX/kk0hgYvdDC6CDAkVmDrdSK50zgHSjj5YH8Ojoru0
KIyliK5O6tRfXuBExCmM7AnZHBlEhCf3tIi/pDfSuTvUXHmB/t0z8bmvTFig2rM2
79vaZI0370JbL46+tW1r2IcKxkK0iu0bmADb1iFGcq44ubhzPdFWESbvzaO0sTbR
OarUvEuk1xs5hWZNIvYD7z4LS8NtIu6FfilafsGEearmQH7CPfn37tFVeyyLxbl0
Mmn1t+hKxVKx+ftjmk3h3fExZ3hx2dGcqo46jDtxVFLLjykVZapWrgUfG4WU8Nz2
N50ZIfOMYuuht2eydv9PzrtLNEe5SbNK+5wicNJhVp1jAsXNpdDSqX3Ez3aMr7px
OXdzB9WcBDFjLI98EN1RFcM/2MexorMy5+1xpLe9OOxYKJCJYZGQE7Kuu+nNhWt6
o/GR5ySDip26cLtK8DQ5uZxEfHPqTsayc92dUeX+3dp8ruGc23d5Z0P17eFh81e4
Ux8PF563FUspgFqpS+VvU9wyrbGKA5dMol0CIQyjIZxDct1XpMSIGuJ/fooTLYY4
jySZK9VFGSLUeQZZPPCSF3F/K00k5c3Ny+m/h2eIqFEiWKg2aSNihNtD78YEhiOO
iL8xnZ8QzlIX+N/uJwdgWnl6O1vnY4UG7mLdN13paNHrdLfI6GIgm7+jLYs2VBXN
w2caUgvVG68JZwGZ2TvA0bGRvYnIQq8t9iGQamLeu8LiF9aXq7LQMRZLTSJ0QKmW
2HU4oXA9AX3tyGYm2wTHKShSxPR7j/WY3W3IkIIA/Ciq9xTYhdX+WgPRpoJ47kuB
z1jeeMR+qW0IBnukE8EK9nRBWinhTWNGpNxyqCswsbzhy5NbBjvQGRw7ykE45W+T
n20URDRHDQfr5jJrRvC3ciOdnBwqu3uuLmRuSD8q2wlVzQP0SsDWtVFISIyeEt2B
gvUgzaDSPhI06eb6LYw1a2uQBZw1N9nfShP0r1h3OktQz9kojUg7Ue1NGs4HIKJg
7qioYN1sL0kQgt+flghVCxcNRas6CcHvwLsGh9ngnaEIPC87Ykhi2qxB6Xt7WveE
0YlAo4wy6aJiZ+/ooDxAItfP7B/HxNT18tR4OQ3xiPq1i+GJ5xxQFdYVyf8bHO9z
ToQgKRylEq7Lwre9x4MQDqGAZsoSVpDkYZKTUmU9JzqDJ8g0S3ruAFIcLTFwENsW
a9/AtLnYG+eGqNQCjPMHT2+iFmdTorX7mvxZM/8NQ4w3+Bf0aA29qBYQW1+3iHxl
e/Vx/k48b2nz/NLlBPHCvsV4K6fkcYawU7Nx6A5B+qn8QhURiGbY/ar2c4/1KAPr
jmg7XTzuTN8IEubHOaY4zn9AJJmgLt0JPF9wvX3CZNtqeV+JOR6sFfTvKvYdi3A5
n5D7e6h73Dt5wZmm/6WXk4CXosoXm8+9C+en3G6/XzHY1pjstvP+P6WtTWMF7a4W
KH9GyHEHcqRR3D0xxIZxlLahOaoNPofp5qDSGVLCTcFzQbvXl0hFOFJBdb4PDeX6
oTsoT3u1ECdEf9AGh8iCUWzPFZf5hCNub2jJjFGTkCHSrCf3P71w0pF0SVrtTSk/
5/ULzIcYINKLCIjd0SUFzDlFtIDmzFxsuJyZOP58bTIhv/7fVRKcMu2HNtSJzFJ1
8BbCDd8j0sKLkgUcdnk2T6ikY2iDsaqkf26Tluoyi5U6XN3EdD08XZy+uFZzsUrS
Fq+plzuGDyuAl94umYk/WXqLNykQkhwD1r+E7gMTqhvIzdRUFbFkwDe5yTP4XW3v
QpGZM+Q8FZewgvfpfI7qWxgDQ3TVUNeGg5w2fZ443mJBM/Ya6jK752J5SkmzAwO/
VXgkMQZ5hdTIX9nI+ZS74c+XMUO0PFbR+zmymOxpvDNNjkN5sZbtdgag6sgnezJJ
urgdsXm2fJO3uFSt3IH17kh1HDFAt76YDKrIzfLn9bpiRy1Cx1ZCkwqtZzVZWfHc
8rnjzWas/i63dPBfD+q2EGsAkzFjRhU+2Wk8BdXNiHDhuHDT1PKNZdoc0UyJ7Lo4
xxspRFxZecYIw2oNpB9vkrCxsPAuAxx1gYCEwa0G5RdINAlj+L+Ic0Kf+MF3anBq
/rXmJ7t3UhgLV7d5RQJ9NRVW8+fuAYrcG9gBUKsetmoKLngMOyw4pmN0bPTBhP/4
KM+LsqhZtumE/9XJIFiAYkV1lYPzlxascXMb6/H72r2Du1HR5c3PsZaJptVxR7ja
1TW1ZVgKMWgLvaqHLcDNK8BLxmPTTINcqAnkXw2yV+ksVlRCYxKydr600ehi+K9T
/N7p2RCcp4DeY9Vj3ycQ/uQavzXfkLqeTt0OWd5KzP/uA9BmuHvM+la77kliHYut
C1wr+bJy8Gy3tECH38kO/EPRKXaSgFhtVKvwbc6byZQBmFrIjLy9MMqdN8buIMDK
5usdAssvZNMCNPLbPTyJQU1RDWNiy4mkPmIamE99BHYYEoevZpW4Gz8nL8I+8Dca
Ts7nARuivHfQgRP18tvC5+iXGOksaz3qHsAiZkX2R4q7eDUyA/ghzVJIx1fRhwO4
P1gWGcUz8qWYLEBWIrPfxN6pdhzurAiy7M9cF4PveoKPye0Uxq7XVAChqQ6r2Yi2
33fxLBffodmLiQutVpJFGk0j/ziYsO6AMPZcMdvVQP3UZzUWGilO5KVl/78AQlwA
E9prcQ/1d7Chc+hFtEmz1p6mBZ9wvOd0j9PzvUpr82Xbq66iUffnSMLkBTb7j+AJ
fQtaFRJfC67XNNcNMbNzblJJPmaEk739h9I5J9cTr5rFLvOg4enEaSpDwzu6xFKu
PqTG9JnnnaM1UZZSU3iwduu6UTNNXX4D9AaZa4sEBMLvMElYXAJQ0TDMTRkZXioz
nBIgKvlQVpThePV/dk+te/xpcMeZOLZdtj8NEfqtbZO2easrX/qKYFmaLJ7lzjG5
/4wh+2jjaRVWe0Ntszrr5RW1uuq/AemPjTT2FtJs2CO8QGQea54ufQMmRiCpZkdw
4pgie57zZLnXadpTtaQ0rLz55EgPcEsXN6dHyCl6YRnyAO7UnbZa9k+uzSfsYWrl
z7gH2fMlzEVXEKQHIc1Z/qTY6bDbKGIA2HXMctAAN7H0aDhMTYZUPj7b9Jh/UFJx
n4dFhYRZ9UbXQrHc0glTC5i3/ehtLYLievtDFoC/5uIt2jhrdV5J90wtAX/q4hm2
3jCkeyqZnCJEBXnl5GhROuw1iRnGe2yGZ0JUT7WUqeIKIqSv/OFeOT6SRQuXQRSM
7k07FxW62dTKCSRtS9tbImr7JexSpvMNmpOgMnICclWoaS33ts6aqsTn6fs8bxyz
a73Wtu/qcCJOqzN5KOe4APr8TFpgpF54EgxLukcTt1LqkZW4MghZSmKY5STRjnlV
gK7RCNNg02h+mlWtOCHZAlr+9f2KSRccPrvRxlg3EjW1IxRpBONVqyv3/HRhkU1i
u4Q71CI3eWBqzaCTtNN/gzR36yy255ZtsZ8QV5kVtyTqoCNsdM+Qkxu6HgRtGi3D
ck1qPYwg+ztPSOqN+ohmEakqPCkfsSeM++1Fnz+lTnvlCgrD86XiIakLGQcgr6yl
YnaMm1ewIoZdbF70rYf3z53VKv+RhvuGMskhPt0Xtd0udpSyiOjn9n6/BJVQf0HO
7DruySxStGiwjE170NLnhuUcQsnbvLp33xW2DHDJ34sxQ4FUY1ketXmC2N8TFquR
bmfaCgPqub+tIJdVMpZjfEHMUIzKuMd3tPRKV6s2SHmSz6yca4AdxfMAdnC2QeA3
KB2YLYP53W7g6HfebJ8t8fekJV+eAXoxdoBh+AsTnbBDBh2l4hL2y0LMa3P05n7l
LRQvZtFFDleptd0hLYrP6hOEEAp+yvD23ckwpoLhZztICrUU5zl5y/oM6YE0N22k
d09nLP/GNyIHxC8dQTH0rgpopSssfPUPziu7hyVcSUcDiU4StaOmJHovzaNCVK4u
ZZtgo94mfUj9Zl6gOFkBb4uhZ6PQ2S8tjrjTCepcJJ3xz90z3AeEXdcGKGh/Ztyf
JKgXmPfBejPf+zqeotUc2JTJlEtsPbEUqBLnn9hY+azzhylXKpyhn3VTrc+58tYU
ugLiCrE6lXg4SwVP5V/MzA4KNJ/X3mOlAIZjKW0I7bTHR0FqA0r5YBkUfCC94aLp
9koA5xkp7/JABZhBV20FJ/9wCcZwTPMXtB3It8BPAiowOX6ZIbDkEADEbYwUuQFm
A8lEpzfrkfAzJLrjWQGEbkzio4xtvggcRd5chSLWMSHSjlNfxdhHcOlo9f7hJ/wV
c61ts/Vo/7wKHoO2xaeEAiUh2C3o+o4pcgSK6+AL/7kOBQM/JEQQNrkpwOSaWKmk
M/ieEfsZ12vcoI/UJPz/o/pZs+RLOJrPv/btsxFBd7vNQuQinLy5tohAHw+JJqiN
Vv5HNfyTMVMBf4MxAQdh3herzzsLSLoaeOb32oo0kJn+RmUhxDaTSilZBEuRG7LD
vwxYPC4rVf2n/XpC3PgXo/AuMWw6kgI8RqaIkLo8WAczAq2YK56UVUH4dH3YR4Pa
3nxFLn6UKCGmPzDcq5s/J2sukoD8qObO0ljgXkQ+8hyCAWX+W0PrHo+d8gXp8D2g
mf9g7EnxCfsTjo7MSupmvFPHzzAmERXVjkdkb6ull4nPPrbVFbaVn9wzhstihI9a
cR06F6ubOJIKlNF+uvwzsBeMJIKMsvAW5woYqsmKa9jVPadeXuI0gpWZUtWgKhkh
RRrNVbT0MPy7mZcCEx8/GwmsqDxGYwVumyt0ZNxZi47Xeho1IgJa40FGqa6QOb0O
Ga+sKI+KSzuPF8OBlV4uJmk3/LMXqrCPXumjmStHJDgCmXL2i3N1+WNMrFN1BNnC
2Lysw0MTYSr+yH6XgoAW+V+4jxrHjmt/uQJmQ2sTT9pax9pullKi/ImQBmc1TxVU
9Hiqovp0wioqr/4sg22WE0ui6eOCyQr8wCtsFYn6qjUCE+eGNojojiwDRZIeDNm0
TZNnia+7Q8o0mVc8x5Gu2xJS/heEHEOlieuqhkWWXQjAFmUNvmCfWab3Dxp89Rwp
fKe679J6CXOzPQUZcw8OumV5kmMYJ6zTfmQeObAKcVgi0PMMCZWB7JTgp1f0xGcy
V0cQBGV99liHoTRyvxQ6544aP3p+riVBQ/tIIZEObvJFUEWxFppxdQ2fn4mvGaF1
/uB9WKtjG2rmMsXME5OHEX4NmZWXdW9+E7QPe6HrfNXNB5E9uDJs8jjItYeSlSOT
w8gmqpzfVMldIlf9tisy0L5x7sGIp7QCUBT7MsxUOBunMCIy63sgGLv7/SQW5rLX
+nGfnhD0sM9kqOi3mUZnrOgw5yu4xgyDdRGB09Y4fYnvTQgWgE2jaKererswgzPa
Xo54b4jNwE5AaDT7Uva9ffT58m8dMoVClJBUdj8xod3+k3tVBPmacEMiwuRQmXSM
r8BYA+tuCTEgrcRQqp0qjgYL3v74QgCHsU7wbWGaaIRpO7jdHAJfN1Jt8+ldfO0c
WZRqpEdgsKMxZU07h/wQaWmH9vlb5TPnkda7P+sy1NG04YjeBPGXMf1kB1tNIy7O
G9t27q2fARc+puSBwlEqw3EeKXy3l7wsGkQb/HYJH3FLFftVaTu05wxNpmE6rNPc
DxkK5OOVccwkS9lQ7XBxktiFfheM5oLFn90n8nwEL1f+NYsUXVypnSPpWNdTxpuq
f/MxXA55riVhWzi5H9tBfIwySoI2mRn9ZzDjQV+fW647uWTbvjmk5CJ5wpnOlbP3
6RV/aLTEe04GfCEBGCx5D7j3lDttNm6EBurvecW3HPXS2F3SXKVHosgaIi5WIVJO
SOtL5a90vqwWaiK84f5TvJDTuoQKRASC6ubLeZcLU7mgL+SotfawmgjBnpTZ+Vfo
blrc2tBLVnfZv+ubiotrc/uSsZbVG90KN5Ogt9hRC7fHdf7wLvtlC6j948oe5x0m
+j97Qpw9rE+hvFV+f92mEx1J6gwGOBYQDsvKuzSUasm9spfObjAEgth9DfgQBY2K
dqItNLlOtYxWl/t99+Tyh1mGD3mdUIfnAN+QDzg5x03BEMU+0WkmjibCrLnu0obN
SL17Ss6A2t3iEZ9HcvszvMXIAlm4/xsMuCkPxS5nT8SLELfEuPnmNrju43+G1PYg
pLT8mnZWsxNmL2VgW8OidVdP44JjylYtNhXr8YjRzqLkydb9t6TuLyZgSXD2LbRO
OXpO+pnJjiraalqIIhcFFfg+9b3FMQ0bVpeXCsjIfIOGc47+KcpTXFhU9KueGpU7
0IA2E1zJRJQUwOpkbCF86Mc8FQl3IcgWjsYW0Hr8LlPfQ9fR/O1zp2fmKrnpugBz
u0FXF0chfV5+JFUFFH9wP5GAEX7vEOPhvj5Z0ZKVaMoua8GQ/SUEhmnazV7GSyiy
Gy64vH4bxvBn//Yi2N5XutLBQvKRARczObaiBwTRx3JVDVPodayex464XTDTKfAu
CkDSj5FUByzmvvPvWcjOu6iYV8j8m9iMBQdJq+oo/WzSlw+yWbq1GYQ6xZJRYknU
PhG6QHPoAId+g997FY5BP3x34ew6xax6Nd4AuHTd58gO8zmMGmmX6b9FVE0OIDV0
GOtEB+ZazjMyRFKHJ4hyZhLkshQx3llfVNZSpkl7O+qL4ddqt11UiSMtqnAcOVuT
vRrpt33hnarbWa89NJYkVa9sBv5ghXYTKC6QbY0suActHSwjbLkOG8ncAs3A/RG8
IrU3ID21IsHsrh68BCbSTaFd23R8xx6kQYhlHqi4vJrmPQNHfI19qXTeyB9oqGGP
SU/T2UmuTGpiXNw+q5QsP9Gl25OdaAP7ar8oNWpVcaoIxGd9TNx8+P2Xp+oBl9It
AAxT3TCs6XOQ+30I2m6cpdlBKY2dFWmZa8iSt7Bvp9Pvs/ZfQDbYvt0YadKenNOz
43OeGlH16iqRH9bseb9ZQur7cUPWeuH92jRL1aaZIXw46sDESbGdU68yclWpRBbP
XwcDexM21hNeNvj9m5dfpSPkjEWnGtQ8s91vHjrXu7lBxrJrLc1F+vNmv5X9++Y0
wg07n/9WrpPVo3G6Ojrv3mef/wKxzpltLUZJj/izpHkPp0OPSB5bApWNYaEzFpEP
ngl4AVjYT4fAFNSjTRNKXsRaXMB4qcxP6oofgeiMMvl7PnLDE3e2SNjNk1GaLWJe
1qojB4dgdrBa9sT2xblZda7TAvRHhkiqmx5DhFgZllE9vStMe19NrIrkkfMMJT0A
/wzBc7MZloAYKV5SkuMqIhMJ6MvBeONpYwd4SHt64O1anhIbASyiz2KVwGFqqtrY
f6B2lQt6k2yBO4pA9MyC+vJduKkpmeC2P8m8L19kSNVA9PaSHYjXIwnRaSuecVXB
RHGaMk5VSR8mIGQq5JS/mp1fW7Iyny0ZTr07gyT2Y6bxL/yddOOmLMYleteies8r
tk/Pq6KSW0n3LtmtNzEMYPDzK+fmbe/md3N5f6BYSimLOl4/iSNJu57KqDKI0ZHd
CXav+N5ZYQ0jO6S9US0fZbg5IoKjxTyjXkjENr7ZIOIjhNesCovwkq9PXbbp9lTP
r4wQwwsMoy6jjaaDL/cfnIf+bDg6T6qynYTWnWeoJH8fuHxKmHQv7Foxl10P9+np
NQTsoQ4zObtdO951bv8IpDETpdAJ5Sh6cxbrCMfBlGvWcW85bMdJu9OJ+qS0hUHF
SarDQOkJv2K7mulFlwNG67+s2VQm97DzRVmWgJtvEOqfW8bXwv60rrMfCDgsYfWX
9o3ZRQqa/HmJZyQfCxVXEG1QwISXJEuWZ5htoBnS5GACpVINrWrePAqayDLu+8jH
QlR20hX5XRpyd2kaHjS96D7rssC+nV/4V4pH3BrEOUSt4CfRhELEK8+LjB8WK8ik
EimU4rQPX1K5sEPtfnQWEVt2rbNCEI1VjTipdAS/dAOWOYDN1mC32+5PsjBGKDkP
b2aCd2J3YGFOLMDhDe8XNGko3lw0oTvoudg8eknZ6tFW2pGcqNxhyelOCvRhxQC3
eBVDUZKT8LydQ/UnqUIxeYs9m26dnqBittQ17Z3MEfBXGVUxr3a6N78xw/bvVmo7
lFMDaOHvgUlTCd8HXgPJ5VcTy+o2bGDBdHEWzc2ZGt5Kq9eOwehygfNpD+S0qHpy
1ndzohc+9R31q7zJkPzzXazLmGQMIvECdQZTZPAK0MfsXQlMSs9Jg7IeKX7/u41t
DJ5IVJKFM0F1KEAQ3d48sgh4mpmF3bDJk5uAtfL2M3FR5X+Ds2eqUhEIsv9tuUnd
OObS234RqEZ+PKR8iaAlaWV0zMT6VY3FuNYDSjvPA6vo5GqJDYojD+JbufgU1XHu
iqPj1ggvi5aKmSzOHxHbOMVdBKyWrzm4PLa0OF71+OACVulHLepu45y54bGhPob2
I4jByEj3BltGBhBu/NSeaojmsZ0t7dIRWAIZic7jT8dgQg5SsfGhI9xDLU6Futdv
nLSvHjg6CVC6CZ5OhLEEJiAVjoOfDOwBLtqyDANODqrbYG+TP4/Z5iHcalbEOFRa
4xctmLxP0qPEhsyt0IWm8tc+nBGVd4h7WG5jZU6MbakD8R99vrmwowAzBly8O0UF
ycbiQpfWKIVv7RekzniKig9MSdu6H86VPMldTayNhy1jcGzDPKvDojanjSfIMwWK
EnG24FbHbGWtzyIyw+Bp0AmOUuYzck8niz0JOgu9o2qwrx19PRnDCCqnmsk8SLnl
i7kuvJ7QtDnErCiKyBfgBuGK3Jtuf4qt14X2XNDc800F9dCFX2UHKXkkc6mxX6JQ
IRmyYPAompdFGRfOPmAp4K5fQe2Ke4ftJ/fy71+JxFI8iZ3LdN7H+RsKFxsEpIEf
NW1INiFg3UJaqBNZY540kiGEWWaxw0/qEELIkRWvaLDpw+ib9n0UwPAvPIHoD82k
wriEwe8DxaMQhL1M5uFHFWNP3TVh9h3i63WVfECXz4l0NTdn/EV88/uyH48nhQgz
5pSKFkIqHrfxs5geK2CMRzLnWSBAV7nGk17aKrgeNFGevZJwykvCpTkmEcB6Bdvu
rGGHs+HHNnxOLlyL/l0JzyxuK1wTp+OdhRGYyKZZBbDAQBGRxlLwDnXD2/0LBg5d
K0hB5R6x7sMJ8D1d2BT8abJuj16kUMG58+dradbVRioIJNtkPQbOM3iZSW8NSNPb
335/f9uY4BdjWJt+QUF6JEH29sbt1FZ1TUYBBf5pkUokkb0CVJQZxBfpyiwj9uAj
BGftifawm47Vu3qXOJrg2db6QPIjAHfOXzZsh2zGOBsSkRZrD+rtsNqMUIiJzdyz
SzmvQnFK+JXpoGrnBIkubpjcDEyykJrGKpNH3RQ3wSl8f+89pKgkkFNN2O7KmcMi
FINMu3LOrf03ZqA9DUzKta5RpsNEB+RC8K/vl0f+Pz3UkDxP5V145CWDoRI6Pbvi
OJyJLKFEkBDce4NM8fquYLt9Hvz1RWF44JAMeLoBR93TNsWBJgv1UDxe19T77Lwz
NQemapN64WO29fY0ZkBmlRTJD1QhVLTRH1WCnRfZ5SkbIiWhGIrkdEWpVxFXsRCP
MElcXsWJWJZiXX5hxZmS+WznfcrnIeq0ZiVKdlg0npckMBZUiA2fxYDj3mTm54DA
tF4PR/1nsHSSHak5nZBOhI/f6UbIItOxa5tGMaayL20JQaIlz6GvT/cWXlqtmVfm
eLxztvyiPg1Ux6oabNgDs3/B9Tn9qxF23Ig3bnwgkFUVqNqtXdhxtvc2x2CgnL7i
6Y5j1fKcF1D1FHdFxULpOPSbrdzbV8R2vHoxhMcCPQ5M4IZ7B7rv7+AZN0THT+Fn
s+EN3zm+LRdCIbryZrZ2tofx9+SP1Fvkp8Ag9pT9uHY8Y72BdtitbcUTGPQ22M32
rLrHFfGGFXQ+TcJz/LMpmQVfunenTu8ner4mDnwlHtOFpSB/XtTmoHbhwdYIVSrz
KcToHOcJTY7tE5E1LSCg6cfzWXPrOf5GAUqCw2jfPdis1hyF5bw01hCHD8R0oYm1
l0zxJPPN7Z4zw7x35vRN0PaMudV52GGFUXLprfEzGlKKlYwzIqtAJmZyA0atDciB
L3QOmGjLR5ZkQUg+hVp9NCNPh8QKs+groceQ9Iy/uSnT+x1E/eE/cCSu2Ba1mQMK
xPY2KjF41XPHDfeJmZKaZ0EwzYibsp3ryHM+RSOWQ2Suio3voZAqpJcUE91plwWD
VaF8T0ZLw9is6IYTEVmvmjBH600DkHyCLyhWqimMj7M4A/Ek6AqdfGvqQYjtCq00
d7Y4WMdDSzjLPm2+v/tSJlLH3Co4/eVxMnRYoDvlxWlZO4JVSK0myQZN7seNbE8m
m9HekR8Zy91HT86SzoaZx9luOG/lbBfJzuuF7Wc2pU+iExaAYBuk6WVc5dL7wEMj
bfPqPqlU8KNF/N68oKWaRGdCtNgKOokB905JzlP/e6jEtXoh05qpla+bEZkX/VWd
nwDLth5XwP6tAs7cbnYGicsoSml9lvURdbLUqnOE2EODG/ZlGkp6mmyvfRFm6cQZ
MAW+6warGsf3H1StBFiVYkIw8JZNUJ/HRbYzHe2jx2AMJ1XO5Zw/F1MazTPULiP9
vcEcUYBLbRBws6bz3ZNODUoZiDY9mOkhkGR6q6rFbdv88nig5clXUWqPTNDRtQHs
/TzpXWOOgMd6ALnqtd5TFnweUm0zcJ0tA0eCYWDtiK/U17H7L0slVP0ZZnPGXbNd
vhxL7KTQpp1C2cJva6At3kaByi53eVtdWhWSXggQKRodB4A0S5SWA6ljb9GjMfCP
9sEe1He3nA27gKK2ujOazPggZN43ZDtCMekLg1W7gPLMKUdgm+/442VkEdtWK7Bp
SqgZ99w7yC8GYYL/n+o6CfZ1Hs45+PJbiExM5y+z5cYD6ciYRwN77PR69nhcCLWZ
z0zcWgbUFBxVftSa5S88NUm3l76/KyAyOfvWsplRgKCW2jGFG7Yi+foGYSRH6IIa
uii/NyBjwX8k6oMgV1/FRUpq/edi84fMLKC3fvE2NkjDYUDL6xQp9QMo4uu2RCJd
e9PxADhFGZjY0mdqeVrIs5nfAMX2tTewobHESoUwFRO1iwTcAgXVvIGCk4khjRcx
CcjZ03iTqkcMcTUrCMpAGnoGzBxXduQ7nqwQb6f1W8iP4uGvquRVCFJ7YcB94czn
fbQLYUIzY5CE+elcx2FDB1kf+1WzWNDTabvkGlQrwTbEOPPPjI+AiYm/+Ry8NWAu
Nth8nzqkJrViOSNsQ0uYfZQgpwPpaafx5yucDJ+nq5AmzjWH4PbekZkaW6JBbiQb
2jm1/iMzHslMc/PCeiNi1Y/6ispqFyduG5UCdsfy+lUnK6vfADuFVp4CXqTgG/Iq
zf4SjjU4QjMJxASQpexqUZ2fwWP2MZODuL8GgB21ITP8LnvdA9/vPpr5XHeGl6f8
5Qnh5Tje2c88AnBgmwlCtBDaRNRGq4puFgxSNc+q37vNeeGW3B4bD9rPERdfNP5n
X1lfvJpgZxwIDPa3SAqFkpjgkrAfUIvKaZeABlhGXIC9PYYr/uXYdl8l4gv22L4R
SblihH3oycv3/SS8EJqMCPA6QJ1EDDne+RUDM7kbB099e83jJhBTj825ucxK9CsY
Omvg1G3ap/7ESyiCWCO5Yc1AuUVsXMX0IlOmq/DeBj2qxS0QInQVQ+x7+kXQJ/G8
G7jolQdqSFtkb/qX16HCJPpe4XRFkJgx2gv16bqMRovwyEDgXNsGXNTrW4ub040v
qSVsiPGO0tK4XmIdF/omocR9GllfgmxqDEq8jeWLUdsYgehgk5881iQn6HS54lQx
KBiWYCNuRo6gAtHxsurwrDyLZgcP/A60eTQpxMKoutUkbN6weQeIymoOrtmXgkbx
/S2plgBGIxDVIFizM+L+bx0CVpAmUKcKaNILzKcQ5DMj+1eTskGigfQamiXbhHEh
8CJpyLct0A7EEdzP691C8kicgvaw2iYr9moBJZXGZ2Jxo4Y8/Fm+2pauinaHk6bI
uH1j5VFVVGKYWjIG8SDDLz3To1I/dv+GqhhCMs1KKqXhuR8prM8My4jXccByKqV1
nQXgBum8EHFeB2PaWGk8l008hIYwLUONazIPBxkA8rcANTunHY1RkSbpgsSrdwTA
EEy4lOuHdAQbtwD949MP+nQNCTZjVgQS7H21v+1wMFa2oixBPgnJHIeiNZ+EHTiO
wwbK0tt/f4uvSmFGe425Jhxfps/rfq74SrRlUxQfQMPp+Y2oWR+PUXtAGpxFf4CC
dbq5a7z67YsdXW9ZJ9+ozjL11WIUkW2bd7vHOa9zFon5W3VHCpSClskHHBlFxD8I
a6YRdM8Ru6TRSPz+tSOA+3ak+RpDoAWGueflPrVC5ue6b5tkeGYXfMMTCxXvhrvP
D+cYDkFADcWvqnThhO+2cAof3ypq6PzmTexFbL5e1QIbBA3nHpsTCCY7HsP7ZTVh
yviXhjFAMOOreeVsnZZtj9aqlOu5kH7nlEgSbamZkcGujt4fXEB6a3KJI+isRzaR
qxleQshNeF3+XVl8itmbWA/XIWgxdiNIa+ivg5U96Psrc9/oCiCebkKds5VJZZXy
s6IEBOXYyGJHjjgFO0MupXhDTNc9hVnMBwq2NP6itSnHy/hSIzcn73AYdV/p53qn
8zWytd+LHq+K0L/0F24Pnj9ptvla+MThPA8Mr5qU5R2hyx4i/xAvYmoON2bXcOJP
70P7cgc4RXjXELvXT3bADnGv6yihOtTWKGrymerVK+WYMC2q10TPvbYV2oLQL33i
/GE0Ib7DOFdDAm0e3pIlC51iZReuKI6yXYg7fZKYsnLw/2KVKZB4qwP1QZXuuqyl
EEG1RI4SBzuiAeSdwUPfIxk9Qvlwja6YrGWBlhnrHhl4alkVVdInGDwXk7BSV3NH
DbV8U45+MxNjLCBTHEa7Qk4RXFNZWjX4GvXJk5ZhBaxaJMqgi66YCWksmM7ILvgr
86x4rEMAUeEk7ywgOwqPlBZEDOnEKzA7ac+sQR5GEsv4NQD+hHYT+kvf8mC9oZau
nK9Qj0d/1HD2P0MnKGs+TeZilkorEu0ZtaJFdG2o8N57SekXLKUi3PmtVfw5bjI/
qsAM+++++2V5Bk2UBqqAK23qts9OIp+L45gw5TXKEa28rKe9ogSPWbAar803xhLg
pmYXQZ7o0T5Cnd+Ak00Ug/qBw54zEmhJ8AUcRu4ruUS0+YOGp+2GTVPuW8qZv0OM
cphDoEg/ApFDsvXJMF5aF0LLkiQ1A9MF8dJr/iiSAWejQOpAUdckx0UIBWjUg1LZ
F8tWzMebElgXgF6eaeL8fugnkoCca0bLBqSIJfP6WdzIrDKg8QlAAdJl0qJm11if
6HUNbgxDaa/UJAIt8WsNqeL1UrPZ1v9/yxm9GgbmfE1tNFtg0q9Nf/mequtMCmpk
Ai4gCsjSH/vhBk0ew2GBbxsBFpystNjdL5cMYuopR7pCW3UA0vnxF74h7bBMORAa
Z6mvRgXOIR2Ft3pzfk8vImJ5ZBBkaFgvjyyLRRwuCfOYIAl+eLDVQBGqCaOBpmS5
RYciycWheA/XimF4BLwX1dJP20fgGLjLRuMfIq/gbWOpB20n5m1wEeHGv65jGxB1
Y9A8t3XHs8TI7TzdTpizYEk2NG56dGkEuug4SjUUfFCz1DzJUXqWlKDbJ9Qs083M
NHElkvYiaADsxbHdNc1dHH3DG34Kv4alUr0Gv3M8EsSwzIizHWXvw+8SOmoH78RX
UXL9Ej6g+wZcOAw1YLSFD9b8ZpLpv8B7Z4Kiu7jfkH2iE/4mkMcSWNiyv0j2s79S
EgAZ1OeWChq2+MYvbIyjqtblFnbTgP/NojSO60OKOHWpNlsby1IPjzsx932wv2rO
FpWApMhtb67GVi1Qxdj/aAX22+qG1BSeGKoWE5B2pI5mPQdRhOhFWl4waGSKQ1K4
IdRuI/TcFan5E1s2BBWDfta1AMAXenBOPppCp5SxcT2PMoNR3W5AneDwiys7jj1k
ggMw1gbQvCp/47/Y6FgwH0nAWr+XC+1A3VjRIg6IKDT3noEH1nb3s7wBcxa50KgU
7nh+SpBHRvfYWHaqyS+DvulixQgx63f2z6i9/9kM31xEsFTUniy92pk1zGynVK1G
4lENEuIT8c52t8I8mbWhfm7tBuPTerOocg/gtD8ePEP/QaSYs2QYSF/DgN/OgXbk
fnQxHbcZKrj48t0MMqJJwiDV1usZnNrIFKrzF+ItpZh6t76q+8I0Gtn2bu3YuUjf
V/2qrVnOvm/Pp3Czra2rVV2QHl/FRR9wWrSWp0AxmbcGvZ0v/m92fijQJ3m3uT3O
hRVA7uTsp+IaIDa2uESxhCcbTHEVySoAXnK7GIpN337VzPzI4qVjs+skrK1TU0RM
TQHQVcfCgWEloUBGUy9xmxplb7tzkRgFKGIN3MDcR4W3IA0IR/IZ7In3KAlApoLA
9m3/T0iTqmmZOgdqq5ZcokJuqCHr5W8qngw4Ph0cUEPwEzEHLcPhvI2wLMDl87FA
ArLqXlxFEpQ2O3tDQcuNZXnLwpjA6RodIGpusPGFXIPFa75ZH66QAAqE1ore1Y5H
Zx6UCOm5HyODZrYsDdnt64ZjoFrTi821yqmYmXHv/Ks09nkEch6apRdwfW7XRgGb
GdORnV3dJ7dvTkglKAggwclOF73TfYvlWJRbqK36mF00AyLuxQRHkYaEgqZZFtZV
O4wEpyPEOoHtvHbshFWnjxGP134KgNuo46Z14e3LCGaVLFj433TOgbW+Lvbqq22W
ieDg1KOjdZs6qBDqY4ZcpluKH0TatEFkkdWMe87wCP12UMI8G8mfh79FYvWfgK/l
h71u1x3qw/33QFXgCO6ARDI9k3E5I4WvmR5X+mmzCLn4mjO1KDJXnmU5CmP02Elx
uSxEv2LdypuAPmuTO/vi+YL8JgG9ITvb8dWU/gnqts2of0FTBq/NVpLTyfBQWqY9
lz7qUXlWeJSqGaHuQxr7jrs//2Pr0LLDhSAVMWJc0wXVbJoOtOj4tUAejXu/PIWN
QwrrZvsMNYNdo5zpgMkyv4sash2jNXDp5PxNuY46924RCO4bC/NohSnpuL3ZsCKE
Zjn+uATFLvIjaB9Zn6PqbJPCbK1bVaZkm+zVXTxYu1GxGjqdmz7ghT8HQ5Q+Qqu2
+7vtAKF2Lk9xHVLijMhk6kkLN5P6nOXNHnK8yK1zuaV/N8ypQ9kM2B7yWGdS2GdR
7eCuSfKes+e/R6fIHhUgSMsSTBQ2IYEjb22GV9dTqXwcgX1iWIiNqir2O23zTIEG
21j/BIYbs7rHzaq0wd49F/DDfegf/vXFtxIQUJqoni2rmvrELVMv9rNQWR/sb1/6
JFZy9jF38x5OzRyanrNI5xxN57BKLA270Syu4sE9iE0soMnYYI8GkPuonWYKJjbg
cd9lvG8B4N9rwl5Kg+1o//NSg7ykh5qYfn16iandMTNgVSqgO6vlK7zCe+8T1KSR
gpWmZBsqB63xAtStgSqk85vGY2GJ5DKCIE2d/KOgd3By3rlAGCb6NuYPTzYwsZNf
YQLVrkeJUMI/en9JjVHMAFqtLwQNkjKAm9UuuQcOHVQMNt4QacAPxX462liMoDR2
7CH3XFy0Yxt7EIFgH/UIOkxqrcUyXh2a25XrcY5PU+aQ4gyJrA+tsZfggn1T7YIM
57pzVI7N9s+GDTMLDCo7bXXYkMASLhlPSSvlc6vxwE5AIuBV5ZjX+nhdf1ouVV8H
HgyDxSMjXPc6S3XKl7YZY9G8T98ns05sIkYNWReGQbSRsWkkhq69PPIpgVGkER6X
/wL6ynEWKb4StMecEivWey75UdlsI39chOdx0G1MpZQr+XRhFAayTPYKGo4kyRbV
B+And4Oweblbpo0PGblXstfOlOv4ZB9nUn9FlcpyEFE+5SC0IuNZ5JvnLJJyoh66
f7sJWOgl3IX5xupUeti4akR2WuD/dZpgD1mfkZvmEV7t1YPxs37ZjoHzA/EhuKIv
CFp0DldtW9360vkpMFQE9KdDTiKZPzU4QYx76KCCSQ2ivFd16r3rIUs9sSBipm72
MnaN8suO53ma+H8iBXHHTH/+9MovXQ1ZgYthzPkNFcR9yOQdkpxGupZmcb9WJOl4
MlieXR4ok330dMQ2DXHIuchOd4ngKJPgxR3J3WqE9U4DF6AE/7C1dxpiom7aHFtl
wH3vXNCmlKFy9fjZy1OP2Azm7zATUvyUEFPgz8mDtLT3XlVw/WerNT6LNN5Kc/MC
ao4WokEdW3yiCyJZ52mwulRiFvNCRn1tNcIPeYwDV2iJ1FP9NPodSbVWc7S/WKgA
MxMl0iKikyj946dVkexixW7ppmhySmyoU79FvnCrRUwm1dwoeWirHoOVs5/bKw2j
e43VPs8pQorsHdtrJirv9FHyqRAQ6MmuMwDambdt18SfFzteHukmC13/vlCEL7UR
y2WzSOH+iChQMWnTJ9LvSX2VBXuB8sXTW/EpfXGlmfRhvZHc4ym7SFlJ8/taszqM
k9Ar/PtI8QrS7p6H6+3Uk/28LTJV22aFTZJMC5/ZII5LmyZdmY3C4gk0vkAEJp7X
vlVF2YOhlu4cr9lN3FtF9PiE4sUqEtHzpS0oeJiNvMGcbMdhK6h4UP0RVOy9UqSC
uPS5015Q81TfxOZgT9HdSqQnYjZiExbCq2OvGXoPRj7TFiKTcIbw0dxLC3Lue0Ye
kjfNcepiyP0bk3+iLXioAUejgpbSrxnxBx7Ssfx2STOqVDDa9+0R+HOlK3DRD2Of
WVbjS00dlRs7UvbuAQBltoukuzPXIiy4JMYxLRUXl8wzrfBLfmMDqvMLwhoxnRQ4
IvrNfjZhz11VH8KkMpfjcaDr5Bru/X7YPZ1jxTeJPFZ9D4u6Zi+0Pk57zW0+wRzd
UORHQkWzrMUoaXEoJxx6xkW74CyImOj/l8Toedz61UFPQ/1wygmkRc4prdx+i5Ek
3Y07LSrylqlxsvHZFVjB5PdzSmSwjHBq2ZfJ/cik/fDUuwbKBVCYc39ly3E5mpRD
yraIE1Pq3M40a35OAhmvrSJsj8H8xaUL2Z3iy4A6eeN86ToEygG8y1xMo8yI8ytJ
1QrXOH6xu1JTo3XL6pTUkvKS7SmXyF9tQauDzsVq4cr+uiEnoIxY/GW9lo8P61st
XBpvbcfRhHRn6n/dOL5KUMJ/H+RzJmU/0juc3w0ITADkmHMGC5ULlpSdNcKlUz18
0UT6mJZjoe1susQ5+EKb2qhdigzMvFBywKD57yOsh/m8r01QXGcH6nekNDD5Mm0o
/n5kx79uQOEZobvYW05BVvs7Dc7+gBaqKwIFIc/sa+T7XHtGbBKS6RalgjsO9r+E
JGaBq11ZOd9j4rq+DfpZMpgjRiwK5gzv1Gl2RMTnhvxcpa2V450yhGFyGA6TgvAR
kpeyP5XE82PwYiucn1B8CMJ9wJ+88kNzoZcgTTaYCsPPuogz9D27Gh0kuOSM07AE
dyfqwI/ui8ezs7WFtAiOxcowCUBRpuOvCmSUr+NnyRSSN8iSukffI7eSKDGABB8H
ZjEClekGiV2ehtsA9chFIPfk7RS0k7LRH/g5+dWNoZIXppBO9g1gwzEah2d6LW8X
bz7v2b0o/iR8jtUk14xTIR0m5KUCNsZZp1XF4RdbiUDmafn9k5OOByIRaGwWWukF
VlktXotLywLCZqx7lE73xzJ7xFXovtGfXJ2AfNC3xY0T6jPoDiNf6AUA8vRvUkXn
6wZGcC/eGsKMiT54kwEyTzCmf7wQ86KYgeyFUxU85AwjE3+AIvhn3ZhFJt7G5UvY
FJVNA+p9GbbCiNHiIZf+OKxXaBjxgIe9Hrw2WfP2zLVIFcvhNcDIQH/CO9Jeh9F4
MeYbLEDzlvwGjdpd2lLrlKSI1unY2gaj9b15JlJTAPuv8SQ0BfCZLkSfFv0kV3iS
2LOOatcRY/UZjO2WmdZtTMn3oPLuUOYeGZdF3YvFvugi9yfUQdftfEdwGeVpsuqQ
JQVEwXDSqD5vmtcfdF/S1GMZ8sECSqxdEvWhz4s8ahnRjzE7b4CB/uAv/s+0I4lb
j3UQd/pz9h8PXUbBFcJ2GfbHdbIzu3eic+/WIsNpQcw2vAvbm46ltJhKqW7KCiDa
q4Bgu8zWKNZQQ+eEJdfYA7UyTrpz0YDDIwl3Yq5BEO8a8twzd3eHEcLc93n6jeRa
hBM9EIdVWCymdg80f4DYmw/6FAocKwPNoxkav3a9Lh75uvWe/Aq/vR5kfUU59A2Q
Wmczzb/XHXjS/z6wEdI93cKeIvRIAtfA1TfWfJdzLmQWUfkOvA7Ve9WrW+Z/m6Mg
o8FucXxwzwvwRUwlx4SBsiRkBEHrklRA1jfgS1ovpXduVhk5+u+Fp6M9zFKCq/kZ
pNyNY9jAhChd/hG5z/zXmxoQjQ5uDINuBQunJlOXD+C7kb3RUez/7up5Uifp+w5+
lUBzrfPq1FZsb8c8ZPQfp8PLxl6RoBitI7w+m+KlDTcCd15PmNtRlgdErnkJFD0S
7EN9cbsEVzdgPBclOXzPYEiNgcRW/QNw1RK6opJtYNJrdowsK7/BXpJQTan8TGIb
BxC9XoVuETe1Fk95pg6Xq/ZKINXrsWDFAdk3/vWXh/88/MSWy4ispm/HOXjPEJu+
0chzcUVcJ65PKT77MKOsV53Pn6U5SMxjZWx0Upjg24I2OIqd9Tk8BTChkRLTtYmR
clhuffDLYBRj1Xj+VTsjbW4jZcrDNFOw40rs3FVet/LS4iFOlvod1+rIcGNNQT9I
6xAVB0VLmjm2Ch+/IemSsvxmaX8QRLoMu8R9j1aBsjQGl5ohFnx4lQ2MGgIigfkE
hSKIwfYZaBiGtzPo4UsYxPZQCfxY2ATcDy+buOWIQRA3MYufyBU9JyvcRTg3uQHs
Ff12TMaw9QNqZ+FtWA0mTc7z4Z/zB5rkhWBmC7OWybB8z6bjQAB5/gW52vvzdFP5
45TpJ3P41ZK4hdqXj6Y58Gvn3SYeaJqqsChvwZhVpl5ow/8tRb/G3rd6VvbtIATN
K2Jf97DlY1M30t0T3qQhU+IeGz3LFjKbUYGHNJhxUj0nH+1oaGfcMIPcQtn+TJ7a
e+bE4PJZ7C2p27Ze1p8rR++NzvY1HVQd7JfqoUgmJslHPzpeCUR2qWU2ekIZ1eYs
YSfk3uGS4wNQH7Tz4zOIOTvltUTGTPD7RNacCdgLYbPj9xvcvX8pGjs/ZTnrtd/3
eHZJUJOFu+0xx+YEfwwUDQkIuQ3MO2xUMDfKRLtR7xpid+Cyn3AA1JrTd0Y3Al9u
U9UdQTg5RzBm+5YF795ZUM2v5OZXYQK5n2g9aeEGrO/cb7I5BvZ9mqTy4GjEZSNG
dw1HPDoYe09E7crSdx2tDr0yvG+6ktIUDdt7IafwCyJiLCR5JOAECP0kydgzypC1
AD5R8hUz4URzQYiTWX2S0+/Z4yyvlk2/TjdMlRbOv6Iqpk1TlDQ8gQJf/LVwL1k7
aM37hECoo4zRZwW1HRitIwYJgBCTmgOw6ITTyygcZob49USfaxW0Givw1HQf26hD
QIJraIafSYrCENAw2BvdS0jag2S6cypnqkZkoKXZ5uVRk5HijarCfdgT7ynQglYe
SxcXABkoMN0wAJefkeP95/IWu9Erlm2XidHW9EVe4GrZeVa/dtgyg8RwU8ihidRM
roki7KpoTfj7bTTq8oT7QazOQ2OlwU/NPM+FEdqPpkwISJTvYLLPaRxmEW58sov/
ykAii2W4RBvqE4jJJOACrE6CVe4/08WgCHs3LCSa9NohXOYqxIBMVznKcj3PnN7a
ZpDscguPIF6Fih8E2R5E3poB26znvMi8wgADdmEYYOa1JrnbRP/yHmB8adMMHF6p
1CSEz0EUoCQj/zOaRQe7lgu2xgbMy3Ro/8orzkl0pW80Yip3ohRVsN1Mq3FNkPfX
EbMgK6Kd2a7PZ8YjAJEJSC2SWPLc0EOwqUa8tAWucNqJyyaXWq6VLpxVuXAboul1
xfH/qhdIqeEPWUVMO8QunfEwNZY7YOaLi2y9rW5v1rd4mYt96Xue1b8qDo2iuwpz
86J4vBYFjhJB+rJjpH/OSwqzF+Kk/nDY7T6r+el0/dmenz/EBd08l/j+WN6Afi4b
ZSHRuCbBx9gCRajkpipzjmmWoBuGVzde6U9PR8T/HSiRmGhwlgnz43QQhIQX6FBD
zz9btOyArF4Hj9QoXO1HXyrXx15Cr/uOtGeDNDsJr4h0E3p7jqsgbZZarwbr2otQ
ltMjSO19oW8CdDWlXvylhqDafaMUlyysQ5JqMPnruzCSmCZdCgTK+kdgJTKSgO5z
ieaxE3GYts3F7uygsXjlD1Ld6FU3hRkDCNkYoCnO2pTJ1WnC+Bkv1y5wAQhQsm9J
ZmvU5aOqHqvleT3QyJJrbnbdo9UJB1E2xUhjaYQ3UduA5kzRwpgMj1OZCi81TSew
sG2F3BhxCtwV+zwaWPnuEc3IyoFdUmoannsfDBNbnyPWn+uF7Cqmg/wT0cpACIk/
eKcLofCSNr+Wq2P2n62nnjWpEXCeYtHCpTD6KkQd84aZZJO8TLQNKvAoe3NWdNF9
a2R6cbgSD5uXhXP5WjSmGaaisbP1JuIS43RIeuYhCYkiLxQLbSyBL/ZKPmKHFDd4
lZs53vrdAnCeIkxqYsUss/3LL2RCrLk4k6G05kMotA5sNUzWiVyevwJ2RkHo2aff
X0efL+XcX4wSXxW3Ye5yhe3mmkFXQWFycu9X8oRgOGWC1Ar6ATPtLWSjGve9euJg
R6MyximaNq2xXAIisbxF03elTOLOB8dyVdzF94FFHVRAS99gQQf4jFSWclcmDMRp
fa3+09/+x/tBcWjzFc++QHSA1XOLKc34LnsYSwz9/kPDinUmLWLkTOVMFxl340R+
XDRKPLDv8diXOwTHdKs6n/0tNfwhJ8BRoShun9CaZG4lhcULPvDNEL5vDglNa/jn
02swgXUXqOqqwHXiK1cx0pG0rT/rAhAT50UMG+qCoSBbEIT3+dSDv31o0br2MzOK
NA7Co0y25LUPBPqJi8Cq9L6rXhdxEnBgjq9UIChHOrtq3ZF7OtBU5rJkeEvhVca8
EGd9FVis2ROiSoGIQgvpqYhKKz+n2cP/nf3cS8KCj9FGjtIY348Af2RxRA8K/EuG
xX+wpAcdj6b6Mti+Tsv/ja1VJnp3x33MtQFyoNlV0ZePc72+bh2woiVV7juHiP9l
hWCkzHldXWRFdyUiPqECGKJF5S0it7C8l5YtEws3I9THjdIfTfpLmt+P986LeLnx
Zq+dNWyVbdgHvOknsWYg0lI70iXUX0T21cI4oKB/qKr6VpbXjWR85/QU0rTawRml
CLedUX5n8wSxhKKYNXx6rS3O81pIR/y45ZKlOLf7JsO18/ZPfma5T0HvWeXgSktb
K6p0tsD17I5eBRCgesNlY/0qhvb4Psez13bQD3gnXLN4VQTwRyFYkY8VVt+d4wmz
DQMkv5xapE9TjaaF8/7skRX8bh44W1PSJ26q/97kNjH98qViCtEpabZmxCF7PxG0
hCNdqI6aPZ6VXZrDVsBOcXuo0oDSkbRsNSpFdXWdnb373M5UUC/4ELLwjUEwXnfo
fioB+JfXJmXaSuGUxMQRbVeKzaBeCJ3nZin53Ysfz7E9+xgXhDphb4kpKy0ZXRuX
u2weKYZGdOpjmYPVNM43mTHft5LfhS5VpJsrnu83OIo9YeRKjZYA4YkGWRRhWPsX
SJ5Ni/rMCJpr7yJ6/pzB/GcNHK5cn8tmpbl14nnAefgKLXOkzvjOzw2rJP2H60Gp
IukJol8ksMVUJ6TwFCJgcnify8p4TDFQMJJpZWIwzeXxt9VdnGHRRdcai9+1Df1w
Eewz+eS30dD8G5Zmxuapn00FoY5IzgN9coAW25WKkUImt6rnVJLq8zi4p6LW7a65
JbnWtaGx2Fai0CJV9g6Hp5gxpBgcg3SGCsbJkd0vSp4wFahxbIi/5ysIBAxxSXVF
wpowWjWbeCg0hDEf1BBL7/Px9XQKwZGEGHLm8f4IfGkfNmU0AWL+88A5Os2sCIA4
qIbBxzKlqLFkSRoCFK/p4uk6EChRDO0wK0VEJhSMfz+FVH7zyXn1uxDfcFGsQKv2
CKorWMU5dKMAjip0b7AJRQOBkipA4zZX53G/ywCSileOy8hfdQZb49P9AQT+x1Sz
Ia4G1tgux0jv9Z9dLRaJzYdD46+q0mYGHulbCXTYmDJ/564qw78AevbYyZ7sQz/J
e6sGAPYQ/yCPGYlai6nlVSTmzyHG0ytq2POOatXZ7kr9/BBrQOLBYEwIiBSbj4f1
ppmtolqhtYUqPAUAt4BAAkuhdqAqeNQHqPE+MD6PG3TN92QRQkI5BSlBQVr8z+07
eQt4aG2cqdRu2+HcZpK0dg2PXUdLVYlr+vieuIkfXSUx8DlZJyc647yuQNmTC3pV
StXf+Y88Pw9LMlKGHJJWrXuPcd1GfX/Dy4vnGw4V171/oTqdELaGz9msOv917uyl
7sqO8bXOy4TuqKFkE+lwwdGntsaSq4UjNqKBNPq6+2VnKNik+tc8aVDCqD4ew7HC
d2Nis+wDrJpqcDWBewyQiSEz15wefY8+SAdMN7x8WPkBBshrQaWMeILCymtIGX0g
ofM4/5uG2CtYYlUOrgn8TlerLW4bxm35ZjVgyxBmnmg3v/1l1ew3rZjFwjE1okHG
yjKWa9xRBVNabK7DGApG2nz3j11kYUdMQneKZxLrpHAw6BT+1J8gssazNIfMOSSY
kWCHBqHauf9kDxP8AhhBZfckflVkrpprTUZoG8ZaK1orb5amb8H8CXvmOteD+4Ls
7MaCsIyeHmEetPTHMgk8wKQdYrZaDMu9f0emQ/GqOqVEPtI639SgZ5+Yxy9JPD1y
tV7imrmFkHQMirPr/4HHmIKh2bC3MjAC5OPK7fsgVc1cMyS6Fcx0i/LBFqs27bNK
1aIYrm6KyNVsiiHegwsrXJPuU82cKHTxSGfmuVbwj+TYzTrWtCMP0rpikbVfZc1h
/CS2ONrXZRcvG2Srufft80HpJavB5/F4epNugzfqJsDTG+MPSQz5Sit1jaUgZpB7
NYDVlmhI/FRVtmaiRxyeLCBkS4qWloYJgds5kIcAGp3kkkGmGJxUBp/ZtONhUcBp
itw2iP5zfFQeK+N4lB71UHVtIeeOjzQ/i0uUrTgbun65y4ekwa4qQArgcBdr4uMt
69rGWIM0bF7/Va1TxKxkXiofpRNwTrWN+93TQfXcRxVz4c7jo2+/j+I/F/5GYNvK
lCnGTeIBgYLUSaKbrgQpHP2OJ1Dj8Y+8zLeghcHg9xl3amcoeabL3LQ33Yz/Va3q
EgQlkjgnOCAKfYgxcuHHIvtgRKDe/4VdSbtVtzfPyfVt5sc2zIFnuqzxcZzK0xnt
M9bAejQ3PTY1bvOiDNxe8n+3021zrZJxKA1rpujf7ASW8Q9VihUvg62h856qgVAJ
hWD7/3ELKndRpnJHkHD8YdNXFfyWuLRaGQ564oQu+lwQv7xgPMlTOSmw+DsEqFOu
Upnfs9HUMWul8EXGJyHeoC+zm6SSmPFBmVGMaQbKLO88toX2H3za/xdXTQCGb25+
mTbWRzPzJXIWfQ94VaOzWCZg0lIMAmYZRK+/+w9kML9fUISvECiEt1wdvWONfTwX
nJpoDFzHP5kVfCOlCQ9Uz/5zadznyZ8t+jTM8A04eJdsybWrESl5A8vLMY/N1eBs
q3rX0rV8CaZbP2zpRCNDfJjm2T9TUkjRzp49fK8MYbWyOK9sXLnvT/V84CwAf3lp
QEbUtRFoDt4kcftwTgMVsCQE89AST2Hc/NW7182DqvkjCN08n7K5uU3l1yYO1HnO
YfvIP6WWkSfhcwzmyvQhuajtO8whmrc58gRRTGnyC6ZiBWMmtlSbd7KclIeLGSiU
OhfyZNLgSq6L4k7C5nEJaCEyztsUWz7nHn4oD0oBGHERwrU7qSk78xafY3JsyLeE
LcQ1r7VY/mMUDTMdkR0AvY/FjTRik/IT2EPb14l8A+wwKBSoUP9ZY1vcel9z9pLz
3sqBREn82bZMWj5Es3V9JnTp951UfsXLWxbVVEJNhcEkJ/QkVPEiU2ORzC89reAp
TFkwbTiSSCzxXjIHKGngB4lVopCUpFtzeFyFJqyRJcPnIwcGYZ4s91mzFqSwU/LO
hnbLpO6m55svkB+Ob8lW3ZAgqgJmD9cxHLMBmEF+CPdhGsjzbdps+N8w55H5SF/h
G5eb+6KzguqVf+q2/Mci47zNp95gZMkKNf+bZgvOxN1Osu2wW3SDPvxTepicFiwm
pWR9SSy5a5nSEc6NPh2VEGVYjWG2epaZEb/NIhaAL4yAmPBaKBI1GgdUDa9PTlPc
Z2q6xhik/t+W2hV4g5G9AuiYWle/MVrwUjF32EDGHiW4/3EGu0vB9kucfxURs50s
N0pXrhBh4MDJVxMhUXm2580TA9+sLjGwHbnqofYKb4mUEJ4MNN/ZNpwbsfocCc0P
SwAZAGWcSelQOeGfe/5soGsqF2KK64S1V2A5EpnzVg0vVgwsaw4/LE1PZ5iixuFw
R+PzPWskr72VWX5UHpSAPeXJhcImrP9b0xsmMQ7w2iFy97/oOJ7EJ2kvZ+8CUePD
sbVggH71s1Kv3prndCdDf2cZ3v53FZRaTLUo7jG+kEp0Mv3Qk+57FtZAYMLRBllq
WIRYnIeJd9SoOUjMrN1kVEFVWUaZxQVvj8YwSMhn9Xo0F1H85dBTKxmLSWc9VtPz
wsz2x70tCjombkc1ZkFKNjIRNoK12tvCasmXczLcsb+YrBCtG3DZfSKnvqySmLaO
RX8cOzD3lOi0PgM5qWruPI3Q9y6TY6DCDsDFjselDCjF782REPtnwdr1Op/SvoOl
S/lskyZ2gUTnVxcFZogIUPLNyhChB74SuVCQfYmahq3XDf4wFGhKzWjXjVK7UE3J
Sv4t3hq6BhP4Ujamxe9jQYSLzlF7iEBVRlbrIjF1iNWrS30z4adStPTmWAsaaJXF
8UHVZddZd5MCHF+B2kFRONnjh1MsuFTbKV3I6xhHeroBoL61/wZ4OQRJ/ruVqlHI
37QaerqNaAP4UZDLflIfZCtqNgJFUMHyc3fnSHRJhN5GSLwq5ViV9eEhoNRnaCmF
k7tZwRY+huBg3WUHvaNy+xtzMz4C/SO1ww6pqIrCTR76LE2Z06FqbADRGgQcFfbo
oX3EoiNWkqtCL8SzwHsABd8b16TQ2uyiRE8Eu/LRO3iiooKfVIJT/Y4gx6R1c1DU
gSoBME5AYfALuPMZIHxmO/5B2oO4PjvHp+6RYuUQz8NfWlvxX+XrR4Mi6TGt6/Ed
i1VlvJWMuHCCAB2qESjOR2RJNjBY0nSSOhzDG6/o2mfXl2xrmLpT6evcpOuIePc8
9e5d9WjXkbkji/ppvJx/oe6Bngmb7sOBrvPJOyAe+wrMsbN0ieLsRbg20RslEbQm
LrMmJlRVLneUWhZf4rqpgm3lvKoUD2Lu6PN9v2qwa4AdhSDl7zH2/B1LSe+VkK/2
x1MXIUvg1VkXHD9/n3I6wtSkueRUW9yJ1yCaaU2VFNZKGJ6MV2ZV0BCOr/nveAah
Rq8/VRy9lVITn7TC4wyadmHjC2togkzIZbh1PCvyx64rvVnImQOhIock+Hw5e9u/
KDdFoDIyBxEMSLqBwhx95yC2o64qwYt3A2Jr81i8EzkVqz6Z2EFURHnAO6Qpzahk
MOXLjapnQeI7NbGO9Xc6TrXGU9OdPXTv567PpnXJUCQgIX1i9PsPtpG2bMuMK7dg
RkZrVYiAkeiygHeplnxTpptqwZLvJ168EsXaoVwHH7jKcAUyyznkImbGiCljTbGx
9g8HnfXkYHPqQ7EyuR6Ok353QIsX2DJpP5VZF9287NAyxQrQCK1OUGgJTUrho9UD
LZNK2Rkfg3IZme+uDB4iHqLE9b8Ka9oaZnb25P9YrAtPMkPpclIdeO+ycPQdG2KU
MbpLjtgQRSMsylxQKZebOotYo8RXnDTH7ETBQrRfMge8+DVATynOeB9UnEi0Ltkm
JIqf+0Hic2eBxyiS8RoQcqKvcTxZHcgHtHTFu1SgK3nE2OfAUOCyXWSpg/2hQxhb
opLLm4UeLZHu7sveMnSp4Z7tzencouxXqP2AZG3skyIrH+f6Sm2Qyetbf5DPLVsN
JSYLl15Ppa+jvWNicFYk4iWVUkUovPIzZr/o/vZecDyXRDNgNcKrZUiO4xADYFOi
dxOP21/7i+Ru4Pv2JfVld8KvCvZGsftSzLRf9VZiffTKydP8VxgBIqE7ZFgQL7g4
KzlGOtMsg6z0OCkr0vGiWuuzcoaAvo+1ynaVaGUnhbXLbfxwbKN1FHIb683/2Qvb
EiLC9dJViqb1AEHvLSPDL0P1jQ3y+r3+CTltubIBFCpjXVsjuTpJBOWEyUZ2xEFX
a2QGDkKBhmfez7rFQTStNV6L4ttFKTIrjO7H546akDChUEPNeUUM0Ls347AroxXY
CRK8DuUeyA3gQzjZU0J1SMHrNIEAgVEgIbU744G9DO6Ux+lBCSPGyEFqK+tbiPSc
1UTLOajf1nV3x/C1OyH1mXIZP50w0BHwVkQalouy3Ln02OZPo9aYzea5CtLOfZpH
spssPRLA8qzbUCLLJIpE8plRhUvmN9X5ZkO1qdn7z1NpyBI5Ul63BM9cRg3RDLCc
EiTIjp/Jm/986+ot8m/kjpvuK0MwSy0DOYM61KLtHPW1B2PeKmfH6vhpy8lSxtgi
ZBWDOjXdah2JYRF1dgEVOT1Znd4hWsnIlaKJ7w+BTYv8DCurPjlUpgn95HCylbcN
GpywSEf41HtmwURYY2lE1bAvvDBg5bscotNvHopEC6lZ7az2H5QOXl6R+fRVj5BJ
a3z8VJKmG5QoLpH1esMJgBdHafEwLanm8oVstKOs7CQz4gUq2t1VGUB3JOrRUwHt
TI310eXSWT8wU/yR6aIXpr4WeE1h6OYGclSgbHN6ag9eqyyiImK2+qZWcdPfuBqs
JRQCOTLC1+zEcu0udRXzER2IFFk1gzTbhapffQ7PW48IXer7Gmy4JgHuqVyN+MwM
cmwb1iSVRp/6VoULl3YwTYwQzs5N/gi2il4wYvb80hguwmp29mfFaPWxthF1rt77
HUC9lDzXa/sRmTtuAG7Fpb0oGx8/wrdzRsdnM584stsV045SaLrJ3UBmjKefAVtJ
TJGGmtruBBrQADD/zr9a4FI8XYZppwvEApn392rcw+OpNUzg0w30JfBz1m/VqIon
+E5Mzce4tVcRtu+gJWgX1jDk2lhJDiOeSC3w/OYL6lknVRNTvRxy2lUzaH1EsDQT
3x7BEFSPB9daQ6gd38nDhC/vQlko9AQirbfjt9ianWMnaGaNNNc3hteQnEoB5HDU
UiRoJrs14DLmDwIxhWUi0he6poklqITNWd/s19tm0Q9blnGnXW2bt7TWyEmAoHNv
LSfaUG76jlf6NuYtJHQxQyRZsTDiUJeO4k2Z3QkEEVIoDN0hKTBwVEwhU4n8XWAW
0q+JLQZgrh6sEIwfucK5Ks2EejNoUUUPPX6WsFgJqvFLRQXgsY+wKKmvtgQRpcsP
eCvJBvQOWY4BCZhzyvuu90b9QSikYYyUn4jQ0NVsEYIXMdshLcGLDHPOJasBt34n
kBxV4p7VwC2w2Ht9MOD3UkViVUoV8e4Z8k7WiXuJh2bUy2GCljcKzpxB4wOqi6/k
WuzhzRy2qAtd1hUXb9Gm3tbY/sYKafypBlY2DRHo3DjTkHUTGehE7U3W6C8KB1BF
U6sQxliqsi+ZydtRlO4PeAGO45eSTxgK0tN4xy9mwoCiO7Rn4KfgknCOTQJN8Ggw
NyScKngXpNoTejWYV+WY8XVBc37v/9XzAcGtR9GGVxIhrd4y/5Nl22xvmSTnqTBP
yPTej13JNqGRMW8D54xEbXiLFmSfr1zLHibXPfeMee4naeBS87/+yoJvH6u9ozcV
1R9YxNNyNJ0x73Ee0GKLK4/pUOQ6uRpaAEyyOGMuCBtwHKCBbBU0YTTfg3DjfGx/
fwcyM6nFLVHIO4RkUcVXgUHYBjVSKXcbpThMBd58W+X2ZuVeBAnavxTFpZ8glush
RF66Jmc/hx8dCiiAAFyJppOvizYFVchoFbnzmGji8R8kk8rYnHaRrudnZPimMyed
s2GVYX8k4GgHUKBGL76vP82n8okyGL7HHEr8zOMpmWnzAWrqv+D9J0ImD5/MmtCV
AuYtNXTWBReX6T6Gs4FfdajPTaz1ps4072fQE4j5XBQ78M+g09mujAdQL2vbMpdd
aFFryVTRlAy3a8sHaADzDFSTU2lB0JDnayMflk7xBgQEk9o7t1i+AYRh+NTDGRbr
wsxSbTmt0TZUoRz2o+zMN6vf1zsauUEYXhSIBs+LyQBsDFz0CdcXCbhLZeUgTH9C
e67wybWyG1xqYeTLYMdVA42L3hhXVZlhAMKuAxtiGZqaS/oa561a7BgidMUWgiOs
suqAJbkq2lX81Z3ep4kdJ5zJpfcB6zSICQbjNtRQhVMQ0o1WwUD0GprDYs6V8bRC
gFpaJcUiK6GPMGxC57QvPCak3luqwFpnNPmLM2TUU9xy0C01G5+ahFyzSIV6+0SM
WaR1Rz5ErYOBSNXE9PBQgXPzosZ/a9VEU7ja73fma/KegBngCsDvMAfQO5YVdWUy
zDco+BAfL6RcEYcQdBTfT67p/+fw2e5Scl4JmQIPzwLY4+MFdoVqYuJ3aixrzDta
LtVqcrBjvvQDcKiPyW5T0PS9dxcD24YrFD6Ba4RHDjtVCaCbh2+DAHUX6GsTjazs
3ek7YaBpVsiHw2RlhoKBv6zkJB/c6RKeW1pB5QlgoIY1qX7x7PYpIb1/INLqH7CO
6k7n7CbPpuxu0OzzyU9Itk3w16uOe8k2j1vjlGfUgyL4Kk0DnoUcYsWVVyRIuByU
5oE4+ywhALpksmoNZuUte9g3PDUAkf2XkEdfi8rAAnA2yJKuOeb3izJrW0SL4KZh
ZC0DwRVZUCX9bfNw9LP+bYg1u2z4DvvRjtgGU/wAOWCY674H9mS6nNKOHW1E2IYA
z0CJizdCEbH9n6qqI6iigaJcpe7fvWH0tX3ROKlL+jfAwS0HhwVwY0UxQid07iM7
Jeg9Nuped0YZW29YxKDAzUHalF1RhC0PIlbWwE3+M6UziactY5GoH6D7kxV+XNW1
bTKJg6aHMFqlSNVBh3p6DysWLoYYPvOw05odTO7q7ZrUi9iqW7bE/lr1HIaDHM8/
mkohlsrvR7EJhTB8eXqilqL7h4cn3SmJJn5mwLEJ4JW3zEpakY+vC0RhFqmWwDTm
KT+YiVJI9sWIOYuWASrNz4DkrLb/VKvbZY4knBnDHt/XDoA/1G3WOdxXqMKPhiRB
x8A8HlnmJwA7D/+antLGBFawLbBSOnVfpe8xyAA2sG0DT1OIC8wy8evYlmAmtiW6
vb3D7hXQfJBJDQVivFmsgqUUxV1ZqiHYWiMZZLp+iKUog8jVw/5J3funsfsALT81
TkNsvQ2aDgad4L7qVHNNNLDAUmHDoKxnQz9w9O07wPlOixbvKFKmOYqicz50K+aZ
QZhdqSkl32yaQM9c1MHZrIl9rtohhlub1XnRK9hkB7JkKwh4udw2yaoHPMUz2uI5
I0eWX2D0ZD4FtxSaZNaGWbLed00wyCAigWsqvf42GmcwE4054Fq2/WuF89TZCmN4
UUAiYusx+c0Gr4qQP3HIyX3fOtmwzGdpVKqCx7eVRZQm0bpwKmMaYOR3myHHmW4p
HCrGeaohfV4WGa3w6ApB7JaN+dfKMOYBjxVvfE5wOsR9EwC7OpvAESavUhGq7eey
V2JW44lbeo6Xp9bVrHickcQDqceI2dEZZMV0zShdXhRKQXaonN8HbM0EVHHGKl0b
ThZTY6J86TKbdPFiFkTbzQTC0CeYbyrlfFPkghExyf6CZVyvHlItMhkxP19c6E1R
u/ubVRAvqwP9huTpjTo3AmcQ/7ntFr7SdPRrU/W8sJvBEjHYvAW8cew3bBys2SPO
HWJ3VpqIWr+n4YyY58oqGs7A8rXAq2RB7kb9jnXvpzf1O5rYZ1yER9px3lr+z4Hw
6IaFu7XJ9CatrfC3mB7qUdC7xTtcJTOpptLSb/BjOeNo8aLewrqhixovi+S0DWpE
ieDydn6Zgy7v4rYguCttUShnwKy7ULgV+56fZoK8njN07crm5khIceroGnGo4v1R
Q1o6m5JRhYuDOiimM3ZYUaDX6s7qEYMlMR4NypUAMpiEPeQNm0HWtu2k98xXl3K2
2mntd2rXI+BJHh5XHDpe9cS+/cS5HwnlTI3+CVhF8TFQCel9ewYzpMhqzIYnQFvk
ERKZaVEfL0NRWl0S8a5ycFLRYOYJ76fDDogUJ1olSEkWZ+6jDZU4Dg5p1nhoPuBn
+Wk44E2GjbfhNy2mEbZLukKhTSvW9+qKCJAhPylT48p1egkczpxbp8P1GrQtObWH
2m1JoiBW3PqBEotxMo4edxObk2XkvsFFJw5gj+QRuru4n5FYkrhtly5A4EwoxFfe
WGt1KvH6M24hEirqM2Yn8Wdxp0tSjKUsD7gv6PUSb74RUW99Yedu26/J9xHr3Elc
F1A56COgP6OCo/NdBtQgKzIsOzgXBLg2TE1Jjn9+deAtFawYfjjpgLtPWhRLgvMt
TtpiFVxNdWQn1KP/OO35+JI8vHgmUqggTRUCWsm4lEhflGB3kAnXSl6EZNBSDHUa
coaU311HlXcU+UdbAaQ5dalHalBBCh0TFtinVgXeQBOMs8S2yxBd7d0Ch7+QO36s
jnO4HJ0hoGuULuF+M/TGTnPwb4Xx4rPdwJxtE3uhif1Cb0VXTbfwptqDKzK4mDc5
NHUdDYQjOb1nezQdH3lwu+prFba9CqTFONl/dZoRgKxb1GCmrPWO3b64B1wdtKWt
C345ncyQAZrYQSPiGXkjua16m4U72lL6g8J6c+LvE+ZwECWNe2UhQoZyj75Xq5RV
lIkFqkk1WX+4/TB1FWEIr+efRkw9lo6SVoZVtG/jN7SBsFh0VkacBYF1cWEnXUCz
CSYY0BG2xAx2DiiAQhMviCXcBN6YAlawE2SEu+Yw9g4E0NMZX7lldhXXKtopGJ7A
6D6rKJ4RSs0lOALEpg/ACjQfqXsdVAP2qluy5SN8PAHZ8RKsE83IgDqikNj/Hnlp
TUn5ScBCfkEOQoPdxZmfAOpEnC+fI4qVhUDUa8EeSGlOHWNdYNa0zRWVRi06JwEy
/X/KF0Uk0XwpOD1gmH5IGasiXV1+lofdJzn5sa0E6i1OnhcBFkDTwHBjh39iTnzV
zgJGaPo8nVWcjOkQKVjM8inGmpbHFUizUqeMhEh2bFoz0QVuIcDvBXXXqq7Sx66L
HpJl2vNZpmSs6brFsv6X+8K6u3LVs5dVcRiTXL2Y3R3+0ck14u7GzFQ6pvZ3J3Zx
RDNzBM2V9sAz5pEJF274KdRO9rY9ejZQsaGj1eIU9qVTshepiUkF7T1u4PZ2ZraI
d//MBb862vWkyfIP5Yma98wzJV7SOu8n1slI42dJjKidTxfVcFhfDXYSWKZ507WO
GuV/tGegOlLJvYFC37g+w2YG6nPM/1BzamFH7eKskG27jl7RmCUTusPYlU/HLGD5
cWExW2O+01az68z7Q7KAl6CJGIYBsyWT8dQ23OHVw/hlx6D/WWGnmbOoKLdnmsdO
JYZy+m7c8TVzHLe0PO+N5FhyQSV3xXR39i7O6Scwa2GL4akswnUVgz29jIcRE5Q4
cmDRopHwc4XyNMJw0m7zLV+0Kk72sZw5omHfzYyQNSEjPjLOYkrIlhLGEGZEoUMU
PMfVal+7I94Z3Tc+UET/O6VePnwjf1oMY43UnwuJlEXDtZeH/cdstAFOJl+6Kjcu
H0xZFtmVtMe8wXNpp1XJpdR7toyu1eKuVT8lSO++CQGR5cy7SsL/w5PCzn8yST+v
dEfXDdZF5YKesF4WuL0YC7tHfPA5zEDymFiwyElwSCQwkdreXFuvll+c174oWHct
QK6GZRH1d340kW2v/EMW+Yps3y0SVA8AkXE8H6+bk/q7aoBYwYxuW9FGS4EyH9+S
aAoBoMIkJGIiyov/UtxOL5L20rx6dGpjB53N5PxIqS9/Zqzt14ksAZAYPTPUJboy
RBtdAbbTPIQJwFdabX78X0fYYKwOUR4RdBAUNA59Qe53G7p/9908oE1OyGlTiyob
Qz6fBBeYg/J0T/DAxWlqGtjuTr9RAsMkksIDCsb8j4aIegle5m4c9QRUxuTwXqWY
P/0CiLvxmbzDbsQtoHDln0pMuf57Jad9LLv41tEd8WkMYTw5+nmTCFHSBqpCKHHt
sTezhXq4i6V2yFdeAC/Kp9aZrbjyVd1bAl5iY5mwm687dnmZQbfrVogBUhvLKrV4
o/jSmB9akvpqa6/NXYsNCRpDjLlXTX8LjdAKfuJ96DwQxhJcUXsFKefW2HOWVKD1
metXFR3yiGFEew5aebhTnUzhTCpkJzmqsN+ORewCP23uJYoW67bzIqhGSz5K5/nz
J9s6M0v9QZPjPl4z6dtX28hGVYSn55uF+5mAIQ8eng1KX/2sw1JRxhAzI16hx7ve
n66DExg3Wk8hxvqZ1A4Kx3nQVyUzB/yJzq/ksyMdskAY5vbl1YT3UmqTm7+69MoC
UKZjb2pizcjdQky/X85IR/TVa/CfJ2TDG7i2gf+q/VeoY+Q3jd7ii4xx8OlhsOqQ
azrhz5DZqonuCeHtkL9nV1JIKo/j6YjyOPzOXavGFmmxfI0U0hRk3x5ZzEcJWroY
3yshXQ7sJFsdBwgS4zSODrxgoswZEbPuBafMlOANpmjma1qn6VJ1lUm1qNGzVFRt
BklgO4LkkO2YFvgClOX6Ps6ub+xxVZxaj34DuyKA2mn1lkfRG5tzXrhSoC7AcEKB
RI4WsS+Sv56pDeM+RYzeMeYNS3ZsawsreNX5YZ3hAolovqcrJQ+hHWv5Eot09JI4
QNt75why+3AFHXBsKRz83TI2EQIM3moirwb2YsjrjZt2FJf5sDnUon1H0TMM+4/b
EnPRdtt+OeIiOHE8HXqDs6ZrdqnlmyOSMI201XlX7CYGujdpHQ2oUDa2pw7jgSu5
e/Y8nbOwRWD/RIIeusUIz/YLsSSuQdreHHvR9WDN5SIXMeyHSPjwuQ6WmhJ1fq7g
LNik9rpQSSnwM0eubDRRDkqCbf6tb4ZfiQeHMg5IauwWKm9oPgj+9StmeHCcqpI4
bxjuE6s9ijK6Hs9HYWT7m6CVRMdRGHXR6RSnToNd8meD7KPmO5JKTRHBrtOG4vqx
tiMHGL6hSAG4Un1chm7vkkzXOKKmQ0/55/bvk0/rh/lzZ94SFWoJSIrtnt6a6Lwh
QCQf54FHkzat+MzVUtZ9EzTdvoc6QNVr1VABMfln0t0eQeu/mxZ/AcSJ+RpqvR9b
y9B42V8LtyT0xjSoT88C92cCUp2nKcUf6G+kobfVwxSaiH5QaKq8ZXSkDAHg4AAu
LLfe8ZqSXgNU/GEW2e0gj6R6P/rhFvkOy7+Uiba4QsNI4sI9xN1Ciw1iRS2ve/x/
nu4Bwlxz6UJEnLDgdWZrdfqL21YS2rB8Bzn1tPPOzUQ2ePtJzUM9y5ZYNIsnG+QF
5sb2sorKvx0FCuvfBPvPKl6jobkIO5Rn8rrkLAPcqPuhW3zwYUqWx6190/jOBwAa
ACQp5bE36CnENOuiQsDkIEyuiSZ0+guiA2SGlh6/Uyd2UBU2UoNjbgPEfsajMbDH
GshAm7iWjfMVt6I1g1kDfIv5zUFX6J6ON+ZuUayT7OXUUX1d7ycfby5nOiC4Z10A
uzs3WiU7UkAGgKW9zU7IS180ndKK194BxhVdw4/LGA4riB7I2H6FBP1hGSU4TxhZ
wr8frcmttsK27LSZFVgXzk83Uyqx0aqzFiByv8UhAZ9naqxkRgD5Ywl+XPPtc79N
7sJowA6XyU5VTOfVRz1YYFMBQcSA/QtuwHxHdI2fg8xrixmedEVxOnjroscp48XJ
9tht5nUKgil0eA65W+AYDmJxN+GpitPckLa4I7eCsq9IG6RDwS+LpdNQq47T0B5L
6y420rOoEiDM4/nF+udid7ItkiGDeBpie3ISaO0qYu2TtmJPc3cBXzlwsfXdsvYd
oZrUbILlCZUd5ff5M+27GgeobfDnUkFZOlp+tVBGkxDZn24/oOvP/YvOSSCc5s8T
VqYT4BYQ7iIEXoPbCCFvCayKolkwm8jWpYs8g8UVgRfdj6fbXemzl85vzXhUH8Ti
YdkRZOXnIOjbFfsoHAWZoVFdjrUOhgNvNsXSYsTelEh71+/d6XWjjL3gRA6P+8g+
xwoLi+CYTH1BdAVqoPgg610b6kp/poY8mDo1NqvWxx0rcOjstX2V5O/4zPc+cjIx
kWa6rM1oesovOst9RoR4I9oMcEi9l2rQgaXlt0AViucak4FmG8EcJdWelK8Rs4Oz
wEXSXKok4/mJpacyfNE7M4I8TDChBtnRzblMw602II1IacEWlK4m0Lz4Yyrxolss
xaFdMBsCZKqV48sNUqJx3h+LbBVkdOvZ0gDp9PkUKHRIsvg1JNuVMMVazzxQqb/K
YWK+eNySHOC49K2M+bw4kXYVWwzg/KiNqMVa4slKQrKq1F5TeK3HIS+j4g2hUXAJ
TG5sdYlhfZEMt33WJbyD49PPZbb08jPX5hlR9S56ASHEcXnXAewzbZeK8WoaiCdR
6aj+TES4mpfFYEMmXzLeHNnK6LfBeC0t1OlqfAZVZvWpkgT0zOsj3RGpHjSkvLmt
eBo+xyu2eUHAa5A0aMtGSLgGLTOjo63CuMlcBsvOX8G+sIj9SJC0SaykS7UXAcaP
c7XZt3T8sn9p29/IZDY4WrbgOZS3od6D1xHRMPXjcLkram14E7RPP42ITw722RQ/
4dIs92btHkAulxUSXDwpP/S0tnjBbp3QXtLAt3GAMvj5EDF3SceACNItoGMozEpj
Esritk6cqkUMNROKMo5xWMeqgjy6hnD6R9YHnOFfUlCTqxSI2DD5y+fzfkB3vlLM
Ph5VxO+a+lTiX7sLKBLxo/xFu2KXZL4zoBnynpymc+gqhnDRFIi+NvPqpFWn/vc2
5SK88izDSbdmsyyBum0tN/lkJ2WCcjcjXuSXOwu+QVBm740xe9p1foeiUykj3EPK
vpuq/EgR5uV/8vquUpPokrRfp6PJ8nUXQuVaVfR5/JgyLJqxER+IlsRzXbBhrqqp
D6yZbvzJWF0xrL6azlbJTpmXCpZIMIOS+YxhUK+joLTMf1+hBBgKd5uYC7T6OXbe
9sYxFeK23yg5x+OS+4GYDO0L+vDC13uomi+NGYT+bNynnHfmONOb+suKt1ryyjlJ
RqGjI0+9n6qAVWVCQjkeF6Q/jKRu9oNFkQlYnn13gvjn5bLKyboK4IW9ap2VcC++
MjHIE24jCgfqa8W917+AwJJGJoXeBqHtgmwHQ/xbfvu6LtQvlaFC0Trf/IuWRw9y
psbUo18/DDZwYrbHA2tjvJRe91rl42TnlTrYMRzGveHzd+zWRmRxtL1HpkjYFBfl
dYWU858ty8eU7rZPGN5h7gwBpw3wKWyTEJGgL1AzbhOFf8qNSOAkpmoPl1pLXIoO
3nA4vCktqatXM3Z6EBACB2KBiBa9s8if76dF/M7EuvuayfPbCi3KTauiBQbJkJLj
xrwG4wckLX0MtsNpfDx7EM7FIFssqFrEnzktAkbpU2h5vDAC2Ozfj7B6H9hoVn/U
BIemDBJv4MOrY1o5Mo4WRRncT094AB+hglWVFU2wMSMmVsJRX7bhAL5IFKleMCZi
nJTNgZnz59OuAtI0ZiHPNbsQPfKNM1dzr0d9tctW5CKWDh4EJ0B/e7AFyHXyXbru
+SIQe5mXr104nHG5p7my8pEEj6Q7Hyyltv5IUBnxYdoy4mm7148qxtANZvZeIpyy
C5jffuXxpqewJVSweQajNtTo1MxfrB2AEnsR+Wpcke/ycH3dKNGojU5Ck8F2nHRc
C4HyeoJfmxdW7PGszsyb+i8DZrpQmTfdc3XLLhPSsHK9L3BVIZ7LCnnIq6htCm+s
NRXYLCQctz7nGYpIhEOMFHsPh4Godzkwe9M7qXmsqRi2w8JB979fFnz+3XvE1MxU
fCCqH6LzWM82bYsPzkGXMWn+9iptF/L/xrZcsKFu5/Gv5rQ6sXuzX1urkZUpFg1z
wMIDSoCAD+J/1Y0iQWST/g3k+PuDbJfHrA+g8rU/yWhP1ltmSBHh1+tzseHd190X
tagOsHgBs/b90gOj6rX2VWET6d/0Mc+XXsKNe37CZm26VIya/IfekoU6ftM9SHw/
w1WPzSZ4zLUjUjNAIvpE9DKsJ+s26YmFPzacqepd9dpl+2i3fTT13aOVIdA8FKvG
I3htlwm98GQkLVytM8MpghnTfpYR/6lsmFhK2wE+r1t9FINCWX+9G/iHy0t0E7a1
0by4YGnqpF42ABUPVCEOJBMnIorEASLdFXvGeaiBnFqb8zmGpDEVu6t8sGNPS0+e
KMMAfPGSTF0FFcl2TfQivtAWUTnXjx8mYOjERCreIKrBstRMsE2tXweiVECKXVIz
1t/fQODyX/L4Grgj5VA5w0DSKg4GlMOePXZ8sBHMfORecmbEWH8ACrLdLGHhwB7p
fraq7TPly2EilOslomWw96orZikNrNlhzWt8eJBkanVWj1WVJsz5EqiSsMuhEYTk
wrpZJVEJbpgZjCwOkxTFbYfCrOuM7IorYtZIZX9xthT4Yn0MVwYkpRoAQd/pZr+O
k/xjsfKGhdgmBVTpd1astFH7TdvRtQBs90PqOPMCZJ7JnmH5KRvmFKAdJ9cJDSls
3SheovU091oiZDPbCI9Gq1+mMSZEEZk+IOS1KV9YgYbcMI+iflNMC8TzBxifojxU
ZL1ZIFmJ6HHNMLfRFl7LbXVM3bUNfuJdR++GnxsUWm5gERIPLbIUaFC541WpCYS2
lUdVvNDTxZCBPFjNJz/vPajob9VH/Whu/DUAJx9XnfKkwg/CLapLCSUP/eL0YF4R
fCORMMatMGc9nV3sb7Qw03VSJbMLYiUWHouQjL630pvoTP0Q1+X2IzvzcCHvtJoy
aZPVkF0+AZRZNwOxCmdBxm8MqZFdlajA5i075hcguGwmWVId65n1RvXj3Ey/qqdr
/Z+3UoSaplIaE366Ow35TfmpQbpbuiqXU027HW3ycl8AnT18mH1ZEapO0KtgJcmu
746oAoU6ueCY1upX+qz4Dk8JXtVhlOIR4rEl3N9upL5BMekH+uC6Tm/5DPAg0vaR
ZgWaqNnMGcPBdLL/OG8Pcmkb+Gdew85LGkFb5amtL0tCI/9ihXG3wZvA7/cRHq89
sFEbiP3/vXmJIYgxjgoYUD5ZuqxhcZBaUc0pTsfuxGaXJLeiYzPD1zGu83D8OV3O
cRfCkPqrM9btZnLz9wn7orQAxcECstCO8r71aFr8NIRSUz8CSkU4WW3Pe0w9uVgy
Ab3DIUTeTBuE5ko9709qiA184ij8W2PrzlsYxGfBqk60+/yARubl0cyuZ0FFi3G4
2tMmkjDMvbWms85aiwnhLhdjZSiKX7mRYQ54Q+VFwXyyjfkSE17ZVquqbbZAAQPc
pAsKkji8MkTDnj0FfUbf3Opc+uWxpxSDFwWXDWtujKrfL9u9hRIR1N84hI0tsahM
3EUvOwnouqLe7XfDE5gqDu49cO96jMW5Focl0SdVWcCFpXm50hoSWlifla5h17aM
PSGmLMSc5G08DwYv4gAstzBXstfiMsjTatgcoJSw+1F/xgG30kSqUnvDhAXOxEkC
G5ocVlYu41DL6fhYeXsi0b2kFbrRI7xm7kjQ47knAhLZQMadUtsvK0ltduwMn6/U
I7FtbHm/eRIpDjpTxIMQl54Oe/TVdQh8x4kD4SV+DTsl+h5VfGTWseOc8eet43g5
+wweKqmIN0RVt+9/jDqlSSa2z6suVMcEF60lH4PXZJ00j+FUxEMlxdfoER5jRGEb
1PsxfIAj1jAxaFWatE8zhAK2q0uE/OSTUrnY3yA1dbN770PHeAGmx6+uN+yms+8t
eW1PdJoRchIL2ewxkPh7W25SwG1t55sqihkWsc++Tixqi0xUyQ4jw3jTYByoj2lB
yVqIjxDSHDiHwQd14yZp2+NQet118hGtqzGp+WW5EXLkr6NjiWEhYjGiJlkj2Q/J
eX0TyFetyOo2xDv8p0XizCwJCsciZzQGbxXn3MZuarn/nG+0Po58W3rdkWrARTd+
fbf4viAmUiqyUxiUPCMkTjXeY1hktHtIgtf/3nWvxMMl9TnWV3RyrWUHD4gyMzh/
CZBndqpcv9PfsFNQemdFJciyIEtjVjgW80hysfALVs0W1AUklpJHHhI0VU95qIg1
6qkqT2uHN1eeGUBf7bQQ2fBTlu+TolksCBX8agUNOvSW1lsaBtLw9dD4t011cDnP
uN5e25R9xw+wnNJuDqWAp5X2/yTl4APAwPZncieVT1wLVtpSccgxj+Wjukug3cjB
JB96ojO7Dih/xjjUYRYkyrN8OmVh3MFJb+JCwQph3totMqi/rId3QoyGDz7+2CQ1
b3zFmjHSJzEy3PjTwm2zwrW4XvVMa50/IwEnQ6eMn2AIXzOv6NuBq6GESpM22ESP
LMYilIHL0CQSnyPo/GqW+N9ig+KXQ92gampObU4EUpZ5fvwyYKtCu6akuC84KRTR
TJCMqWlELlFzdYQ61F65/FX7FOVqdIqqmD1qfyhfVHxNYadZcUgeDo+pICrEUnfa
/Mq24hknbenHJ2nzFZ++pdV9y4R2aNeDIv9Xi4H8UQoZz2h8H3aTxEDYIxwpK8BM
x+fcC7Ll3bwbRPVp8MAFc00iugsq8VVtoJCuF9GEu0iK2OnYcusWud5ZbujrBCrr
Y/EgXdLglFluhubLxiycXNQs8rbQ2diMGeHEDvnfnTJIuqETRiePnq08LkCWICSF
UTBqDG3hU1OQcBIFxeu3fAEMjGCJDl+45Ut5ZA1wro6gJa1036sUn/ep2OGtHRme
Hu77t8jsENpn3dQD3Kswn1+f0ovth6I5B6E1rIVugzlO/NEwVdNJ4APiv8iH86RZ
u09uBsAL864iWM912kTc2xG7+cKx7cXyBWZ9JJSNjhDex8YJK6YmZUiJFtUws7EY
C0P5aXLNsU9CqocamE+J9kNK50qireounRarYdN7/mMDFDKIIosFv4w7PhM/tiUa
/0ipW0f5oZiL4rOfzOxFF7n4IepUHmHU+N4iCdsjybGN/UjD7RI9Sbe1atLcwAyd
jxfN0G70Q8K8IR8vJkTcNAejEoDa2hpSIJmt86uRXsUwEEAufMy/lHjTDe5BFTB0
zjsMINau+mgtxM+4g7wPGpBO6UvHHtGwusyc86O9tsuwvxPQnb33wtSVZBUnqyiI
bRhrd0YSv0cWdDKNeoYQTAWPsrVQQv/ib+xlNF1CNTsQvMCCzo+Zpv/ZYcju0Lee
OY+CTWqWxuyiIhPKNSYCb1xOV8j9Tgap83lVQH33uUX/bAMjOYW1V4iEDzhis+n7
xT+Z4MPl+w4q/5x4HNvhGoAi6MoI829h8sJCK2KUYjylZZc4AQlVsNQKE05nkTha
CsFK/3ZlvNIUigWPk+FdCPWUWwlqRiRCXPvHU6scuc/kAxIMNGGbxMSNlnDSXkXs
9QA1sxOl1sGbO6DnMq0mw/LFzVZgxKcWP65sgXTaO20Fv4bJO2RTjIm1w2/knTtB
E99OgRyKT5+0ASSNCsF9RIl8rcNN9cqJNa5VlwxbFZP3mbP66Dag4geT+sljnKYj
BO3hg3EVGluXORnBaMxuNFIFsKZzUZVvF0WdiUVtPMFFAqtM6HlXCxFsRjq46Zmg
d3LO6Xdc1wshiQi5Gd2Mc/bqysICF7lV6dy2R0zwy2r+H6uiFyakWwVyMvsKSL2j
yo86jKRSF5iBQJ3RDMxmPUqF1jekTKQIXaj9ICk4dYZBBKngB/f0vfRLfoJWMOXG
o2RIWllRi8LtEZzuwRR1WzxRAumwr/uLtfcvcumWXJZ7/pdbuXIjNv5/eIQdTbAf
coMrpV9MgLgS3gYSDWXpFTJtSj/lDRIw0VeK4TUdPZH64w86GzVVasXIUkznT/xo
mcGM6QqOFO3aIuvQwc5EmT26dBG2CnE6RWbUNMf7UGZ/93n5+oTGRQxhv3gyO8Ev
amL1gvIk8F1wcNhDvVZbmn2sdgpp8M2gtwNPK/aDuhX8vXhkfBjYTb9djPmeFl+f
M5H+XtowQqIpJVJo7kHSMtlA1mF76T4FWQF2kbiCOi+QuuidXmNeo1NR5vsPtb6K
LANU4iwRlUpCwpRpdwPDZ5vXKeRB+qmwmOjqYGhasgEIivrk+6EOtD9Kk8mGifFj
k9nGqLkpI1QOwqVyYiLikrbVd4z8G1plUxmxe8okIpmFBENkhOHmN4uFYvS+Syzo
A4dvfJiyhdklEnpjsmNNnfzshblDeTvAu1v5WEAqXp9zP+rHLIqVWA3HgmkFOSGt
6wWGstUXJCPJSXGS2ZU+Yyl26koCdczCaUJTFG9UhKyw+TpuQB/Gxvak6r3vnL33
HdXNB2sabxjUb1OekQBcaBdTqFGHv3yBtS7ffMjUAsK7YAi0Ucn1OZZzY7Fvq3wC
yrS9KZHVeDz7NbMCbuLJgJfaf8cISNyYZdoO0HqSWs/s6dDE2axFYrlVOBsCk6nf
Tj8FbkYmWNQWn8EHRAVVDRfOein+V0pSWtk+bV/5yk0+glQTd+eZ7ACd5NvOV7ZI
mUevDT38Ciqb5DBxJBG/tqPqlxw1hKcRG7yCWvKnFbeYpYBWPcReUe+kPjuOXHFF
bm3bA12tTUVrCrWkcIzD1eVL3/Kzqownt1uUKrI87e/+ZZeCpBDYz9Ng9ssydWXx
oheLN2c5lyjJalX+vrAwdVfH2PWaIcnpVPd73IvCatX53Y5I2ld4BqKSwS2uCGoR
TvqOWREW9SqBwXi1CV0OjHCDaC+Hlw+lCBv229tEwmEhTKtlTvVDD/zP+HdRE9RP
MZ+j11jhEmhiks/dhcBoXbJjUv/oq7OYeCdnf6Nc/5BwUKXjQnyWfhCQltCZbIaP
n03q9iujLYuyHjHqzjyja6YL+a/6cqGmauVlwu9SKm6yxPKloFfDRMcWMqlc7XZv
Q01Nal8Pqg6T+Y+5r5ENvQD0Kym5Gx2tmt67kRyEZvfX5517Q1cXtWnLI37kmi7E
ebwiTeKMVpUyP2sOm7LKqclxH/XWb998G8P7YucXiWL7IZtAhFfeUC3UUsubU1Zt
iidhnqWgBvCQhg81kTskvRvlYTX5DWqikjKcbBr1v1a/KPJ6HjAs94koGYSbDLgV
RcWBsXV6lm0JExrhiXuS16CDowd9loABtHMHQi539ciDabSF4ifI40XiavFxav1q
LP0Lb7lhgQprdvkzoRES+8EHLY0PFkKHh/hej2G5zSMe0MJrw4vz2tOG7oJihFC0
Y1Fv7xCY/gL4cWYRsp2vz0tTGldiwjDgJoUuYHTh/V5waiwz98MYaCVsNd8OUi9j
GIArH4f/BkujirHc38gid0CAxOWSnvdYZ2tHtRQcJq2km4d8rlNHDFpkhmlXboWA
BqMrmDNh4suSvC1Ni8Hfe4ACpK0ew4nks27iwwAAmZAkTBwrxXkg7PaUwOsxbovs
5zP1U+McDOr+qjfyat9RBqEKiHNTMKNo73oOuo5HWC5cPYieQ+KJsSSNn+VhLTlM
kDhhGBJhTWB2IKYZOhm78HjmEErXS2eUV6Oz3hukrMMk72dMqP883XYXNRSS7Dot
UybLN66IzsFoDgOnWmLcdFgsyfqZhXIwMBW3oLLaFYtNlyw6kwT3et2MbyrSix9R
HJoubHex67dXYFq7CSaA/bFP9VhErhx4FjDpGXA3pdcRhEQvhhQrOrNQe8/XrGve
zxFt7LrT73vWJWya0FT8GUiY1G7mrAmeAIQttmgLat3MrAk7Xx14Kah1O91drTT5
MdbKMNZOgHFgc+smjQc7Ph2n3e8IU3I+T4wNeVdHliLokMlLcKsKo2tyXVKHh2fO
ZVdy0vGkXBA+x/s+rNTzlwvZZO4rjwNwlt/22xL/jWhgaQyTSVsQ77LxvBV8f1P7
FkDEk5W/be8P1rVTwFI50XjkUVRywPcHkyUbg7cKh8C7rozhHRxBC8qXAo2chqR+
RX0Isy2fE9yyJ6iWK73u4SmZwXQFEgaNlR9di2VT+v+pQ3+8qY7YjXdD0fXcHM7E
/txjR6dPA+A8QiFi5cifa3c02/UMNFneNybsqHwTHbznSY3+3l4aRCS/2mfWdOb+
F2Ca9AZDM8xhyoAW3e/V3sMK4dk1FpMrhh2SxGukpfbL9zyuUGyb6OI/aDLwZRHs
wBVcXa43XkW3y7OgjGYEyP+CiEZLtK3WGfZETKstlkXly4MguASSTc6KteCgf3GL
6FFUR63AEbGux5OYBuVAncZP38eRpr3ouGbHiDymZhooCYrN2X0TFuk48NUPRZ7C
VmKU70ATea2pdvSfM61L1YAe28rzcMXoLTdTiz+1diFRX948Jnc8U5ArK4JM2R1+
VmJnb8213pxUekhRDz/rutUdXfcQjlJkVXYatcrJYf1bgEqBBPjUVZHFdfzPf3yI
u88CB4FezmLGUlUp++Tg2iCzufpcoP64xtw/KBLCPIgNejwpvoPIQk6MakShYWoR
48q3UUehqhdW8b8jlEVd3md8W+bk8DZChx0ZthkkcWTvgTOOP2/rBpuHJjFnw9eE
Kh1CneBgX5sdEHFl6qGmlbrAwVoFvOYSAlmj2WF5bEj6h4nD6+qlzU4BOCbWI9Uq
0Uy4he9xNfDnLVSo8ZbV1tluPDgojrIHwOtIgHt9Ygkghhj0/P3VuqlHkPNmkuis
pcKVB7cOZSHYZk104bP6YRTrdXdeB2zBsGddSTlIoTLBfplFJtYS3UvnyXi/XKaf
+ucLDZVOAkx4QXuF8uxg8oaM3IfPUIGfnoJ0dCVCqwVGiJ9d7JvIvVVTV+z6lPzp
L++Eb6jWk6LB19l5B0H2L+S7viPse/3D8+bFqYLSqxZxkqjL6+dvljarT71dMGMw
sIndgOs9dwYekp65TESGz/8H0doy+wX68GObirYqx403rGbyCHJb/dlQA1nO51Jt
L+Jaj1ozc7HL0RYKnosekigD1urOKt3TTGx0xWuN0bkhw4nIStyZS2yyqlJplZht
QJ6jOcPu3RLkOTuMSJYIx5xp9eA3+qSFuJdsnO9ZWGN0wih4prq0Itzy9CNI71cf
T/NPHfbBxdE6QISVlxeA6fwkW652Xa4C9ebY4xWh45D0FfkupkAUFj7DkRtUdSwa
P6DEBIfeBNYHBCNNetd/8db4UpmOxRM5egYGkw39oMTJiNzvcQYEDfRBlx9XgENc
KUVXak1ZKXKDep3E9mxN/Jf9mpQKJwqUOsRNOq+anwVvtPqsPL9vMFQ2+JK5Tebt
PLXwnaxfkspBvgS/voDX/0dyC1cykw0Yt70F4spInl/JaRF4cp/iQJiox1RPeNiQ
oMYnvKXj+0+ccqDae3RajNCuu+eEsYYmIdZejih6eU3ooiVgPua+K7nq/Lin0Num
k+KX+vGcQ97AkjMRiFedKS3muvr7Ev0pZezD/hvXovVShPDjFan8iEJm9dM2fha4
oNjzb2QFvb2PXzYYRMhMacF28g6Ho3TXG0U2f50dsZ9fzebjw7v+dtBkEvxFJooA
ef30cul+jFf4uKH+46jWiArfa3L1ZJO7wDPtnPwVD/S+/bfZLICNSsvdhnQM50IY
jI+jjax1I8820oF1CX4BfxZBkpaELXurcidx2IacH+kX9xt5Nj/oEf7h0HV8eF8/
Y0IXNWkhrdwsz0BAr3xOF4XZ2M28p8uooCNeNk2DG9O2/DYnh5AEBJdeOzURdkRz
FbHCdFLvMU/rfLJZ1lP2ONeiLzY61P3NdaTnsDy2HApgv1zKCA36D2b+oVtI3u9w
8K22/ijCHveNQoLIYIc3Iqf8TCmEFtonDyRYoZ+MbwgXszJmbOHQ6R9aGgiJGgcB
dBxMD0pOwywwUgjq9CJn9niLoeFA+vhFf+9FDUHW74ouPa1k28lXl+4+M/pPasga
19KEt+HDEifAmQkqBmgjZlvXoQL0NHQ3SgCR1kH/uQqn7z5LWqs5CnkNY6GcprJZ
dUXYIm+sQgW/D8cwMGJS9WoG+uXCiPRkZj1yPGIt1xdLLnHcLRhv0ufwsyliH4QN
Q1ZbU3zuJ7hhywFykCRWhiXCFhVbQkh62pyMHqlXKZXgazKtMcSlLCHTyXliDn1P
Cl2QdC2s6iset4UnkJF42Eu7JFFb67SCUETwUI3TQkxkuDvXFpEQBXg8EGsnr4Sa
AE6LGHpPDpVqSRs+E69K5xbPMa9jCBt3zODBhrAOOSvUDVeh0OHkwLMKpMq+Q9yx
+cKkwm3cL+X4rfskA9usYMaqefCQbYPM8KV0e1NELF03z7q/lKwRhDP4TlTcB1GW
YRAywvRnWm3AbYmNWFcL6EbMdEKAw7LLcRFtbqI7XbsRJGI50e0Sqb0r/h0QJ+3u
L9IoPxCuVbZhxtFxCmOxZ3dMEWY4gP/zSAR2gHe+PiN41g359V9pOBhpli6i67DS
1r9QRiFKgH59S5daTJ9iL99/zesENPrYsDSJCWjmQ+b5vbB36XLkqS04FAdtpf5i
CEFISm0FKqS+SCzriSLE/QWedRJxxcM8fUJOUSgqB2506TQ0m6CpeJ3XgHuUK0FT
BG1742sAkkWVA2vd0ujF1q0l87Myp1sDGaDoDGJNj9MVfVbeIHaWLgNxOGuHxvMS
/8uF2lpruljX//+zETwD/8xk7LsIvEPEQZDfDqgkmqtzGgTuE2QJN8Cjh38F6xuz
D8DXycy7c/9ifF9i/Ho+n22E7NZoTQiZ5FjeeM9EDsmm+bxoVs019XCKNzGynH6d
gHEPY/bNDg3X+0zyllrEeYNEEBjeEwld4DfbzvbdF82FAvhHBsiqpSqGN6cDt2kU
WfoDPIILNUkUxBEKia70Lif8deISxcWEavjsw5CrkNQm5tFoUFuYBBCztijkc0dw
8eAk07yIJWB6ttZt7Xf6qB7GzU/9gphlBujlIztKgmIdDag/2pqwkvXAfQAhAN4s
n0t8IVsShf+u93CGDwJ984Edv37lmnli6FN8OSvoW3tbR9jj0rJnAslGkTtMy2kb
VJIs3iNcQ1KEJWgjYxM7L2QomiYh7wHs9vGtETXKJUGyVwcaIe6P6gl6vs4qhPnK
5aMfZHPzSfk3dobn1AD6yW5osL8fn/KzpizbKJ34O9zXcfx4Ex8tHoNdFMcFGYI9
0/mzpocJJThWmCmGS484OOcZ9MAdz+F6FNS5CJ5bxa+hn/cXMVYXRl0e39l5Ra50
mbMdNvoJbPzs5z4Gqg8KFzeJAJfwM3U0NugCkYq5TGPJ252cZYAJ9NEU6PUNNIMG
sT/Q+Z4vcxXlFNwMTETvr04IbgRHoS286n24mnDIsgXrfZkz8mIvWE0XdpLMOoYh
7OeyXtke/ud9j21Kid5MOvUdpuwAVStWuzFEhdKGBEC3xH5T4ErI5KN1Le2Mp/EU
NnPIlXblxfaL7v007VxWxE+gPcG84RgbVDszDiM6bckRaSx4OTEY1BqiMigT3Scu
ocqj14tEBvY5Te8CXSZFRiNvP5icItINRfEutIjw/On90Hk96/7Van0Tqjz2lAvh
MntJWn2x9AdPQvwi3vDMJRoibIrzGOkTBC7s/iza2Uh/0qRhsxJZWW35/6Kyunoz
Qx+xQjVCtYnKJJMm7g6fGw==
`pragma protect end_protected
