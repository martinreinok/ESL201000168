// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
UnV6cpxk+lxqAUTrLNw8o/+KONFbWeqqwJqtPsj2VtE2wjYwuSUVvmb4v/L/3yDK
cS8OPlSp8B8b6sOaNIWPr/wlWFDONg11e/TURxQyZKHrYoe4nV1HeCyxvWbQiGuA
NHeCPgaqk2CHGRw8feElCpGjlXs1a04iN/nczDPGyygM8yfNBKCAfg==
//pragma protect end_key_block
//pragma protect digest_block
n9pyEm0FIBFW8p3N0yHdmdjbdMA=
//pragma protect end_digest_block
//pragma protect data_block
lUaigEx4E4IWVCACFCUS5BueAZBeSk0Fcqtl5HkJin1ejz4ct+pLgq7aV2VR8Nk9
3XTDizAX747YYc92RMC8J1jMz6oi7CskfIixwhTAo68/t6IEjMqXzo8SNWz+m6UB
gMp8dzUHy4WJA0D9CoLbb3D1Mfs44SotDgTsHpHymcVkGOFzWfeVaADULHQ79Sw4
lrDVUdiCXGupRT6S0fUSy/YL9gqWqcmpe7mkrtLflARJ3DCAlsOT3a+pgjDOFQE6
YeQv16gGioFXoOD+sNyLn0wDw/0XRaqgkUWU+tMgMBANp+xE1uef7/imGQM/Oah0
6jqmVri8Q4EI8py2Wqb8YR9QUCtuiVX4n1C4I/GcH0jpGY73jPuubqqKx+Y/fLZ5
0fmBkjMWQZ0N3qfl1qr5qqlJV2Oxj3XWBZ/eCRSZzDc16cUFHk3MnP48VZeEJWEH
mwtX7AMiA0CF8oUlJv6piCz1EGhyNIlEdymSCeENYGxHCpeTRWB0wcJVuVoXzTcb
/360eSFK3nqfheg1NBTby6aV9pOIDbaqtgaqSadhu1fpra2ctFpk1hvy3CHTqaew
je/6IG40j3CunbhEwWzmxTwmybab7DdbrRd0T1VhdRwjtulDwGsP0F+O6g+Gecwy
kgy36oJpm86ejexn+BY3KVISyK6/WWYssIP0wnrUVchDL85b/EjrbR+jE3tnch2i
GuLDPj9YFaUVA0yObCK/1CeDEZMqj2KeWBmGGQyEr5aKyz0AZGv444fh21/Xl2Kh
/uCBEpDdL3lYYCX2RDZWko9LXcRzI3AljGFxT3bG18k+2dViMMxkVTVMyBx/Du7b
gSZHdXZriFg+uXrECiioIi20L3A+hffSlfbqk7O7zlhL8qVVwdMbacNRfyZsDG2g
+hWT33WyxdOw6RiRTmhVLVB4httWY67YGqo7XNS9aGFEBWFFccskaE3NVxZqIo/9
eVho4TxxLYsKGfjkSRvQlGIiM6s3zu3z4P6S5PxsYoHogh8AtI7+nWAnCVOtRLYO
d7NHLHR3kZBl+zW0EDP+y8NU80y+gp+yXW0r7GTJeMBA/NjzkIOuiRlXJ/9UrcpT
2cYeVp3OZ+ZkQgpVzNzafJZA/ATzG6ux3dpQhj8MaY38JI2XxQSmKbOB4ydU8WrO
lv/AAZlyTIdHolfqqY4bu1HG4RAQfZDHDAp0TUpnuWviuEZcXDrw0jQbeCs39W72
A6SfLzhn3I5WPjEigIBfBvobnbDJiU2xqdK27ChM8aRNCIewz9CzHXz0gk9c3d+o
AnfpFjr6H+n3VBBiXWK6a1NQxis9Swn7JriCcxYvOVx6PAZKXm/0RTzP3VrPmv6X
UorKdUyX7v91XE4+GOLqGaPohYcNiHSgTBCTdicK6C/ACWpQ9MvPJh3Gs0rALfXC
NWqrI6ADGl1Bafb9iCT+NKU5Qn8U9AUr+tOsN2azDGq3UZHyhqxJNDmGiMgxCJRc
NhbQGz22muBWVHCTYyd7v9BKJzPUJaG0qxuaRbY8PjD58qZTAkAEnGOcayaXQsKL
3eDxTwIETXeP8gsDPatui5uEFQUbzLPmg7COpeMj1ngWG2LFdOAm5ufhqkqhk057
tA1MQmZFzQsXYNVSuMwJ9kglCYbKN7FVmIqhNVAv7BnBiPydXPqrgPx6XEZsSnum
AqeZBPG7A6Jd+32mLUej1XvbpeOHdSQnegLT+rvxw8F0FWyXqIgcfcXdCKEEulxn
ouY4BSVThSdYu7BpDMu3yImYwZreY4IqC0xV0V7n9IuzqPralJA8mOUD7twqOFDk
Ei2EaG5mymvPlFah7i+yIq8YpoB45D7Ge/JaffgiM9XD2BVELzv6zmVs+JoeCxvP
2f3kczhszzt1Bxrh5thhmUVYGCJovEJJeOS26xdwN/JEIkrFhKsXgSki/AvPkU4l
aTDSUPGku3Y1NeDLD4R5e3AfgDLxxWdiZ91XLc6ss/z6BRwIHuTNVE0l7Ou4kpVn
eZtsS4tC1XKghSVuNCvub6dG5LGXZA66dA0MoJrrW4PaMNbzhnSHUpTQvstdntq1
wDqKUxt/Mgq/werdXi94DKvjFy4jLVUagncGEuqflS3xDhfElaIEaxiIJjX5C2uX
r1fIiTm61Y7NhO92lahT3LMyY+6mJNk+WSxEWtkAJCvrVTYghHpqvoMcxJD50K+o
kRJ/2pMzUP+t9TC0yoR+szSdw+mrkn1a+nO/+GxuPp8/WklWWP4fNfm+8BIECeky
ejUhekzzt+5sTZDVuQyRGUVGm0KEwWNgzHw8V6etNyXCGCKh7hC3Tea2CrWBVWoq
PMJliVxHmX2n9Zj2APaxQdo6LYBYWgUTNB45JPEDOFbcbwO5Qo5Eq8EOhrW+1Liu
3V77iNJjt59MiFPFWMX4DZq256zfjCewi/4GxEXQ+Ee/NR74yvfSy/SEHLHAszI9
3bTfL30b4OVhmnLWp8FOmaM2g5N4aaGaaNy3ujsXKGInBUFCPHYPoOnpW+lnb6if
zqEoSCGIkL/SDX9tyh74gz0+FflE+tqpzrfRGFDWEouO5jfWCAQCX0QkfyTriUo6
05fLKLyp5DnXf53mSbfyx3BQSc/dlbCxm88zUnShUVRgusJS3d8Odptj9gW5NFpS
tmNe7XEH29kuYz/ctfY8BPoMkMG9fVKPZ9jn2r2vR9tavrFREfr4sRFk758NFXP/
7vI8NR+uSNUI8dG9MD7zG8P3yCmCnVla5jmNA7dhCNZ3G0Srrw22Zjx4GV0QXzX8
2ixtgi/ACUHx4a+KANcAEaOmj5gIuvt/MH4BEHfEpep35wR+9UYeNKWV2O9MVTv4
3X04WR06ld1Pj1bd889IopPNG13z0778d3JykO2GhM/1x3EPFZfxvPmjZLrH8Fiz
5bPLvDsA1JNlbj7sM3Ggnl03CCGL0OfdFf4HyybbBDEryhCYCm04e2fh0kfJ5udo
HTD/GFziAf715VKABH83i1nFSLpTpoErPMXdE6LiqoDb0pLhN/t4J+Qb+Bv2lScz
3kEm9zOfHxxsYOoJITBEmyx33TL5hR4gZFUcvCDzM+LnBQGERc4L7Pp4epA75++z
OpuMD4NYUC02Yxzdrn27DJqLLDe3gIasCPDA0Osyc9ehCWWHzfoFku5EMf4ZNQQx
XMOUzse8A51zkRoMnmiaMCEFzXmPYxttnUSuESGoLXH4HYeFqOCGrjTObEiIUdGG
l67GArh24zYdb3rss55s8QZiJ08H0fIWSiANGvfCbSPx3t5R2DTNVnNvoBXM6/7Z
KTlc2lpAjvSJRr8uSzrSJT3+zKrUc0Jjqv335XWcfiO8aUMwIX0RpeS+eU7w+lXc
gCmh9Z5fna86F+My5ewSAg5qtnYzIIwa9rM1Ar9Xtu9UcQJVTMCbZysnXHn2FUNE
rttrYhbEcFMzT7flXJ9QRvjyAjFg6L2OU+kTjpFom4ZfeP1YR9RtuMfK+Glpi2vt
2SyB+AdcnORP2dlxkReC0Q+5g7s27aYuktl3Za6rygkobU2kXI2lSaIoNex5xwkb
BD8RYnRNzhI+TGTbzFOMv2lfuP+co+UprPLaWKk5fA1xBzn9vhlb8+zvvyZEpOoZ
v0h8Q5J47jVeKet0FDYbLRLX49ecn/flt4wFyXEIrBtldO85qV23VBg3Zw7+bXTm
3j+iegTwjQoKDkLPQ7e4jmMmndVBaiYRYhCtZVqnKehA7DF+5xWPCSnuVtgSCQkv
R47ASPuuk6iGdLKDrWToQMylJ6jxIqIFswm6ROj8Z1BHneYX9MM953g6YnNPhBfn
XHV8UczHs54DIvINo8pa7nDkKFimbfZRwgKu26yVK14+MHIgopjblQu1q6q+Z8DR
l4VU44OnNAuxrqfcBIt9fu3Ro7oe+5+UoNQ5zCt4wKAH8mekAFLcwVNzYokYB0YE
yR4aReSMSIwrBUgkytmoDSMmDVWyER13VO4dsUeyuXfPHJ7g2pnNKrttbRQIVsvg
seJozJlnmqPZ8cKAA3XzjdIzWIMYzahRvZmfJjItGzzmUlc9RZbpHqyvbBnutJQJ
RLJr8IgJlrjsRB+nP7Hthd9L5KLqsfO0aIO0KradE1m795uecyf/UwVSJVMkY91i
fiqU+Na/BeU8UnMbxqmNJYsTV6d+WZXQlLZDtRbQHpaYUrceZil9pT4pTknDHcIG
rzJWZAk9PKQsW7bijipCcvY9W7wiPlXpMBVNcTyiUCkrxSFDMgflq9WXrHgXQHPf
T5g47juk5m6w/gPWHmLsnt59AYix3VMh/iCxs1UuHMpVJdaWjVfJiT0txgoKxdQt
GT+FKqx6Vxa6XNjoR18kGJ8tjhXaTK2F4dB8kWuy0vwAgQ/qFLkVS1jv0VZRCXOk
6A+LqGxuOqhFF9SzW/IlJ/buCh4Te0bTA6Za0Jz+xlz5EJx6X9Z61Ez1aRlbdEUu
jc/suBDq3u4HKMn8ecwJnV85PB1XJ9MngPldV4ktBThMvH5AiumVvenOA83964RP
0PA0beUNWduvLFC5oIOrOw01Yu3yN1usyjuinjiREPQDrTbMSIKJf5Gw33ZGaCJO
3hEGHL11//eXX/fhiC9uBve1NkWyCSViCm8jhXFFfQoN5JeIIjuCT7yKgjehEbqY
j7mSotTeKHC+fHjFOLiwFFZGRBT7Z/PKb8H7knMD8EQQvjlHimVOhNDtrgybOii5
b2syGiJ8w+OJkUKneWcE5HRx5B0XEfmFSl62z5B1BIgvj2yEw0p3k4nOtT6T9LZ7
1xaL5VbyWqGDqCLouJ1TyFtqSSQnfTUXyXRD1/CSZKt7opvRkO8cm74W3rgDiudq
YgMcy2Atyc5lGDoHw32NLjAkClETuEU3QSpQcuC/j8lEfNnniJ9CsUaLWHXurnmf
L1mwZyKF48Z2jv6fqi1Ma6s04eVtxNvgInbQOBHvl12uKafuDQLmIjkZa09jdmNe
xn47afGeUKmakTIsM0evGYWIA3Bt1VxLX3dAMA6a/7rNhrkjP1IcuFhfgXa/WQk7
0VWCaFqGa27mL9Og2TKChOSG6s3Q6AE9VpxT0uzoBXZIAui4rOO4QzOt/od4T7Ba
ydjmwuZVDFtTngKIfRNT5pUCNC+QRVNSjo0+qXxvpEnMFW083nkFkua9OdtcABC0
Ek0udSA18/EE8FaTIu5vLC3HC9iiYuJrjkPTXAkWDJcDIM/7bSmAdVfb+UxPtbWQ
8Ztfx/0ACGYIv3bbtPwpGnduZLw7n8Ts1YnrLZoSEiEClqySd6WZ1Z6t/fIMutAP
H2LU7LeXcFEeYsSPIIgYxNzFX2V79g2D2GP8KnEMn1SBBpxzcdwtB3wsjSI6EHhQ
D0nrPiIQihTFHdqNVMakNqRbUQeBmjs1pP1VSxp7P65eFZQUYWu6S5J7QcvU3huO
kJHpZALHFQxbR1Y9sAv1bUmfnstzqDj2DhLe4FUQ7I/EG024RjSIIzHLxLKjVaxn
iTPC++m0fyxmycxv7L7o/dN5REig028AJk8cbf/u1RwPuIIvb2nJ3ZyIgXZPv3gO
cELw7WIqXgKDMhnJjISGLCyyTXIee3AnM7SOM+FwpMe0kYqg0b4yUrldfN/q26/k
m+2SGeQrJ9oSMV/EV1a7WY67oJ8q+2OkdYMQPeyVentblJ7vF6EXoEkEbiEvwhMq
SXz65mFqLII6oXtsAvMiArdV0Y1pU762tPNOYEoi7/dQeNj0BS/Jp5FfzwDQ0vCU
DECEAb5o8ZuBdDDBYW/1G9lzpfkc7AiyBNu4XlUGqvtGN/QhuRc5TCqtRCHw9MYu
BPK8Lol4LfzgNgRKms3kKfHpT4xcthsmSd98kvtNjQluKR4hACy+M21tRbKqLQSn
CNd3sSNcVygvV/qQ4t9kdFNy2GsgsEJw3W5CE/TsU3sgLJFWA3X59JCVChMD+C2F
/e6zDf3Y0b4r+jMrO02xT0Dcc+xpTBsDNhsrTzfToficjNqBon34r/cVXBBwOfgu
hnUMmsAt63KD5GTqN+SnXHQPKDcb4hlp2sF9XH8+TAFzyh51Gr42cgjji1yiiFs5
EhAYNajbN3gDVY52zsho4eZkMwTrPK3YE1shUqyQxMv2EeJE8i/PkdjQwp8cz+Uv
R2znon26isWJMofKieYheDIXbXsquBcIgIrob+tHzHbRdjl3kZBwKg8lz/6mZ5Oi
TI4l0L8fT3BE/oIyQumLdqxQh4ndpa4Wg3ypVfljO55M2LNdNLbAb/2XyQB0t7Yh
Xtn+B44XadytuSxBgnh8tJAulNg7jMGlOH5D/YY8Oet6ZobmHEOzWzbdQG227v6Q
6KrJqFTH8j9L18irj75Ilf9vaYHNwK4CvSNKjAyGuVp1Lbs2GKN54N9SheMxITpg
62GKCEgmoRhJUSGDS22OxlhER9g0tWqY0wbXZebf0dQaTDDrS47IAS47dqlT83Tj
Ikvd8LvJmMhTmuQCF4s3Mh8VzrRgll0m40ChggMSSqxryZj4zo1AW9AJLUPu3CZ+
J2eZctCwr+5Jr2Zy3q/T7vdxDLFlOPbI44NGnnUrQNv0bcaKE/3U8l/BTQfU57IB
vvpBlERhEQPBS8wnS5ccyE4UGDkhMGCPYuFHGaNW3goS8pFsiWR8GW+xL25ofKw+
JQinIjXrW9ZilZa9UBVFMOI6gcs/nCgAV+4qjCTnB6ePU43U/7vpztBG6bEa3paY
prgnvIquFk7WxNKaFbk2LjYPtzTJroS6OZGsmE+RgZml/YIVv9vPP6SLga9wY/WS
ResYd6fnJsJwokt0Li4eueTew3RArlQwgyrZdU0b5jVKpIdMP0nCh2Msc+pmWokJ
SAxB2DWUzd4C1LWe9gDCWXGbqS2DWCAPMAUGPqYQkQb+7Wrk4+qHiRWtLUd2Nw4j
/wBMVw+m2UCMHuT1LGkmt9aRxVFfomVJgHhNXXSuddvOj2ZCuHwwrYoo5OMAT2Ay
17y/SAvscpstmhJOo49bmHgq9l/wfkymL2VluRKuNl/e7Grf0pjrY3DsLUCGe+U+
oZDR2oI6Xbm25VL0G/4qot+FqzaOmKgamcFbFXTLLOz+Um7DY0M+FXd/Zbfrs9oq
SfKvP1WLukpspF1m1If94sp+1LYKkS0Cj2BIe7XhcUROvdrX5OMupJTTOI6JLTqD
8MOpAOkIXC5kO6uP8+cD72DLQpJec11IVdAfDBkPRonuWYgIM8ycpTNeJEA/6ITo
awBL+L/V5CynvpBOKC9WpIwAOZpK5RSthjaCOPuXheIvguKJBweUouJ88mM+8+Wv
x7IwwSh0wwd6CgX2zBNnxwy3q173r5Ya2k+PAWjfS0yUAPzREnaCezj6J7TPtKHW
E+gEZzrPXKsK4QF53EMC5E/uQdDRCR28sHoS31+ZCJ88pWMZrMjrwHJMmkv7YKY6
V8wPM3eJOaQERXqgUuNAxrSvrYLL+yPnh/CN0et+7Sxs54/JrYJdWOUE78P2wVaM
vesmdjmIn/gq84smF4eOiQpZcYhNhP4xvI350LLrvTrmUC3H/V0w/Wd34KDMY/CY
A4jmS9dmO1QAVb3kbLQY+AFRpjV0bc1cdfnk/LuuNDSZolffpMTXIA81eK/n9qGN
2aq1JH1cir7AwzJ0PczfXE6DWInrg8Zmw8rsfyd0K5P4ZDuLKe/g/YE8TZ1yQFcv
Ln88Zi1F+/seu3mxD73sy4wawE/dqjwp1MLL7X8HRSpNQczvAF32d77pgHT019e4
CqypZLbfI0Aev5vvWS5qyH2dQ8Gn+sQ5phaqRwFqqW7oheXsRyHvZL8Dc3q5WnHe
pCBXszUp8xBCXP7QNMvlLLr/dbaJGTQH3UNlGeLlU6AuruzM2QwYzFuHP2eT0OoU
oiGapnEkneOITF0GezU689F37Knq7zES5/OCgKQZawiauqHx7FU244rGirNh38gZ
xp8rYdeHfFkGmSRgeZw8qKrOvdI94X30S6CHcqfJmRK/HficjbNVnwA0lh17COOd
RIYDWC5je4/8Uyhk9mDfLeppsEDlKIx6ixhTUh6gvQUvGzgtbEpaq4LG8rn620Eq
AdFzkwc10TLfWBke8ElsZdS12e6ypmueycMQcOYMdOE2yCU2Olu0YUBZ0w/uhrYD
z5rikCVDYwuEX/ionzsLcYMvPyxKDvtkLV0mGUlOn9orMQksRcV3UuKKhE6UTtog
E0RdxurnMw5Uh9eSiCjxLdx0akJO0qF1g/gZzszm9x/2lCJ2YhM0nVB26PYloTmc
DJ/g2Jr9GSe09xbPLC+ntg5meVuSSyL8ChRaW1BhZ+QViyI0ym3sqHXXL37c4mgN
irqZYEp46UKk/jGBwvrak5kU2tp7OLtpvv5sDz4sNFO7QNF/NBMnGcop6bTDzgtB
NL6bMbKbvelVMQJkLduErdDwkkNPRiCRwBR81ksjL9WpL78gHw0pPeD7cntKgPl6
8+Z8bWWTwgISM7zKe70FEolICUL5mD6mSbpWgzRv2sWjPzVoKI6Is+NUy9rwYu3r
tFG46LGJUSKW2v7DI0x0ot1Um/tT7LGD3sIRUxdi3iKJDrvJcVC0ZSjXsN2Etiqq
Oo4QiF5uGMbFeKS18tFp3tkuch4eO8Zs9MYeDvArQwEgYMxSokJS4q4j1Vn0KMnC
00q4LVsrGxU2RajzYR1dKniePZF3WlRUP8UUG9PRTDMOn2gMIHJ741TLKtGQJGM4
FzrWGjnKURv+AfuDiTRfwSwtKQ7UZZMokT3mrfJMSWJHGArMvJB3DROKOk1OePAS
G4jHey25kcKB1k57VXZYoNjGIsxfpR2q8Opm1STR6uG8Vvjc0Y2EdCD5txF/gggi
m5mkL7Hot3Uy0giQ2+L0a0lkiCms6pyjUvn7k9MhvxLbLhArH9o/p3DQ5fKFXqty
jHGWbLNXOHsU43+uLp6Eu0dbESWfA+hh9dO6hfb5Frgl2goHfvyHAzS0v3vBD6CU
t24P7Pfs3yQMjXwv/rby6s1qomWOLeaG24UBRkrSBR6Ixlfy/GJ5fANImPoH1CxU
92WNwxziEFCFiGZhOMSERenkOiIYku3GxCcEikOeVxeCS2kDa6bWXygnczXWG/xm
biQGG9WjujbGAa+mezuipLvVT+8tbSpibNMXCVOy3LhKwDOih35Di83fSPHKlT7g
vZ847vcw8goua5HxZBGl+hy/mHv3i5KQxspHSkFukAh9nCzKkbQa+L5ZGSLqyXnS
lxPsqAHGB+SsE2/fiv2zhBJKtNSfk6a2TLaeKn5AXexumQK4JgGvT3r95SlgO/Zh
u0VXpUxEYrdqGwVk1bxsvl6iVMhbeloqpi9nck+Vsu96zmNDT6p7js9PhxnoO+Q2
5yR6q4eqFks//HxQaeNjYaWNk9l/DFGRUTeyIg86EHogBWNs8EP5YBAtiEem6aZG
d4wJGO4NowYVtBB8HUT2WJnzBP68wHOGnGVnsWpFfDiD4DxDlL9WSbpQvYEQabE7
khz9a/xbGZmvzhQwrRLrdCGqI1HHuPkGSYOXajuFrbxf4IU18CyyTTWc5LaAdA6K
g1b9KK0pTgM16Yl3CqlrK0zEflPTGRsqymUTS6eBQEx+DIiPRzlE7YyogeLefceB
yD4yvntuVrzPs7MJSO0z28uEO9OKhKpBOFrGs6kuQuxiO126uVbevvUIDC4eQZWm
A3XcP3SM5Jg0ANINc2SlvIE5FjSlF2Wc509+ecp3TOVOrDk7zKrPsAZwBKpzVIf9
jqBxagmaIz+ERKCer24jM/iZ+48RASFWeyEsVYrX6EF8M0W2T8ndM5vIEjor0DIW
ZFOAMD5tIICriKfPuLcMbx2RQltdvBEJpd/xjkRRsE06lpmQtYZANqJkCCkNNz2V
LUngRG1zVYSsimLV3arG6iEhmFrHbjqS2GECI0yeiTFGh6bwEvTGxIsLYiiBztoK
WG+qEDtvQyG89Ex83KPDYJDg/7kGK023RNyZtJAVuVlK5jEFO/2WR++GkVbr7/e2
APWowcnlqaNpXjTYo/h9tndMydCslmx/e7GOQ5JksqOxs6RwfTKBrtdEHeccNuNj
4CVbM7J3mln4OxzNWfHx0M2GJ+aJLxRiwMkDau45bFykdr5rxOYQ9ewqsc1UUGKf
9XGcMjCCjjdBOHKBswa7C2OM8QSYxz9cRQmtVoglcFUOu/rFmATPyX6xxvT3M+e2
4oroE7b1oPbAsbET7wAFynV2uqQfCNgCSOnm5apXq9bm7hcd+NTftUPWZVtUPeJ3
UU+0TUSR4NmGcAAgfVNJMu0TUnEgqzw4M+qfUUEF4VEYbF/jUPplz+9BsUrp0MDQ
ORQ2Jx8eunoQr1k91Vr5bbHZ+3EFW2bKP0OoaxqXEtRkGOMOZdmqoP5zfxROXlfy
uA7bJwStfdtLaNJwGmsHeodg8t0C6yRgFFhEItj/RimBHmHYmGtZyGCdwQlogjH/
likT1oh60zRGEWwLukw+g0D5RoP7Bq3J3f2ek+mS3N5IhuODxHRo/qsNWwDAKIQm
YgZYARXCOa02BSBkylK7fQGSdapBD11Yv2aoC3+mY/ppT+ylEwqXMul7HHpBUqAi
GT1hsBnpj74EC6ZYIS8QC5zheQVi5fkwpuDbFdyzciCqpTe16LL6fude+LGkIs2G
GF4KrM7VSU2O6bCAwjPw4bxL1cvMNtI8MWmAqVMN1Ysq6JmVHyaFPOHDabOOnldb
FppkW2XeTxUAyOwhrjVrtzKVUTdQbmP8pK17BJVQmde+F9qZA550k2r60RRjPteS
zEZv4UKRNIzFFRV2Xv2OkqhoWfU7SRIIPszvPHO1t1KwoQNhq2aTw9fEd2KXoik1
BSRBk8MgwMcwqyl7KLLyG7H346UCf0cKL3gWQFoVlLV7IHQk2mm8+apbR/Lvrkb8
zBkoAARLnpBgYH9YxIpPwIPaffMYDL/O1HowhIrliXWr+MBuankQJeDHgAYE0uwo
4Cp5G447fC+4shbPYWHx8WCb3g4oHOqX7KogbBEnqkllO0l7pZG+ViMdD0O4lHSx
6dLh0kfAOVyxAq/tgSgtyGoY7t94snOjy4N9JPCUGFpyHJKsvVobKA55rptJaH4T
pgkPkACmtLb5hYWS3GjHqNBQu4Y98WlnUY4W+MZYuqH2rtwYCerBG1HYtFEKay7z
0Hi6c1FkjCrvDCGPTLTxKO9T8a6hweUCIOTKBJS3pgnmGRaFuhykeBnusR5j+KDG
Br+kknuIpKGPvcjK+aycjEhs12yE1yPYldLmOFu3qaxlT2oGKTm/lxrdBSDoklsY
wZWUQIVqKzw3uPGHwmGOxlhhbtNwrEm6oWKjwBC5c3yZHPh+WhGOAG0nrd5RsJDl
Gfm1zBmIVzDjHmZF75P5LxtZcSsZ7Jgk5WtLHuqxmk0gjMQoMD1YTVrEZFnc9M2s
BXdR9VzKeNUWUyk5yOtL5dbezIwFJBviRMpc5I3sTxChU406qdA0I5NQRDEx6L3g
07zuuDJz7HbRU+wwbt8e968OCSuybocGXi762IF8P0Ak56NXT/FAIC2ivOkoqotC
hKjoJpGUnhAPp5Rr9BM9zKF0qtZlMcz9q1KflyM+rOTNh1XsutOshuCL+tIR2205
dZ/4i0+oXO5gWANk5yJFMyP8USnQzKAosT5gBxR85qLAGYRpFiRC+FFI1U5Y98UG
lpnqgGNNC25eUNIgxUT1pnqoa6UbfbPH9OdULfNMjW2dLNpNz4cmuYegWIHdLllQ
SqqP6eXqth4u7zvqnKVP/rwMlrhqZkJwWwdj5xFYSKvDmvJqY9LmZcH0Vcr+mQOE
NOxAQNAaMxAFvhf8GWPpwyGSEF/gsjG5dVVcfAe5fDEwr/WHvupcHypBjpabEd00
ZidgGWNz3NxFBojNAJFGBTns7BNddq8A65QkEnriV2273KyydsQapqst6ohevxCf
p5yaFJgjzLYswlwbFoXZOg91BVxwP6fKLT1SL6NDDiFhIv/A07PfEC1fc6tNQCRj
B3PrU7pc3eID8x821yEV/mewQyY+tl7+sjMfFW3I1nfAXECWUSh7Zc1ewzXiindC
/gtXaFMCKt6Qwq3xExV7EThvxw2MBQvZI7Q3AoYiIWuM/9ooEzuoRhao58mktJhb
M6jxl5gwCX4m7QjR7ZsqHQ+T0kM1GeekovwjLjUw5XkH3IVJvLYKq+i9OHWiPzOd
gntUgFee4JoFSXFbseAhPWSAdBosVelFxYne5DRuB3rnd38+b+IVddjF588pK3Qb
hbueWtKXgj6JLQ7taOd8xQZoolffyNB6mmY4OsZ0+ZKEg9D+gv450tH7kvuxoHt0
fxu7iz5b7Gw9t0d/yMD9u0Rm2WkPhijh8NwOy/9btmkRx3FlnyjeyxpERdtSE0uV
P+m6vHK+9ZkT5tH5XQzo7iy+TlOuJcF6hsINib1b4AVmk4BvMFg8pRjoyzkC+NAW
W4Gq5PZsp94zhB7Hfg+545OIOacXOgMB6OSan5vYaRjZilS9V008ubpxg9mX66ox
AD6tLkZL6nis7gqCxaYQdlPo1O4pK5C8X9NpzcAv9MSevV0mHNpBccezaLgzsxHW
beokxO5/yWS18n5+jXkIQBkZjmK2TmiZSywAMeNoJ8Bopcn3mvDb5CuYR/D7zuFi
PLCxOz/5oWzULCzh9uFC5rTvkHatC35Oa60XXcqkYuVFUQR8GDSmLuUJbIV5nAxm
GfhkRm6sItq7tub7wUspRVAazjaOix3ANAxKw2A+RB4QRV/eGDpgp4BZko23ayc7
C2JxNMQ5bS0yTRfTdw0mlQDFhJIDgj2bGeGvWbf6nABxkGFo4QmZblk0UzLnsVC2
PtLrOmSkFdaMlaG3ssqoTOQS/f1ZGVUIbrANAE3DNbVt0IeF8qgmuuth0bviSNfk
XYosV4Arz7Ua2JOYGRtshAXVaTr26kzd9hhzvm56cy9/zSdaKD93wh/WETPTxCsV
BMmUwwEBtKFgowzOIBzOgpB8Oco+f0xMZuhn+b3cD0tqafQPhnCzqU4cPuts5rcm
jwcv96G/WU1Mp+uu8tXrQSXaDHk0J9ze6u5iBinRNpsjwDTFxSCYaQau/AjGbfMb
wPw51zpzNTsPcAKqxH7BC7GB3BKGZdcMjR5tDHrNk3a6LVzrJM5/gJuOHZQx0kLI
+pDsolR+1Y99USeEx5I4cRyJTxgeyQTwCBa8DADhw1U9PGZFlvavdzKk0QIdX5g5
85mNF9qONcJC7XpFtxHto4SeWFX2k9AjQEutiTmTCPnKwOa2cU2OhGiw7RvPql3V
ZJXZDSGECmgTRjO5nPQwkdrG612tnJI+5OsxgVUFSKl78vaBVpgIQRNEtlz2WY5+
efgbXo10B7eRPMZG69I4ndrg6ROiHfRBimVglNsAXpMvjOpCQKJiVDONZmj8ES6H
vnPo26OrufI0M/q0rVBtrI63oZr2PcydfsEuQ+cbZXMrbGmUekTvf7HuYehJDt02
/DHPD0jz+hbnheCLpOGjWs1UWo54q7uNI+UEOw6J6bPnze8NNuPv4QHp8hV/3f3L
PGnVAd2H3oR/LjzTKtpBD46spH0NCvhD43L8tP6w5+SSIemg+m/bmYeKLJbuWy/l
9VFR2BJieeF4x8Q8Yice+IJPHm7xCMjVCWPVt6JvIm8+npYSuLmCDOha2tqGRe8h
qiKPSbySo0F7fdVTLkNobVFp3lazPJR80zBoVNt/P6n1pEbf9OKrRsOO/PO0QRwz
TLiQxF3FrQObOfD7BQO1bH0/0fjvMuL4F2RLlhhE6cEmSKnXMhfDTOi7hqNf60hu
DDwLg9+kfKuPa6Sa+FhjHS2pfV3tkO8PS8vjcFr2d8GQZMrcM4PeHqO+n9qFVEOb
xyE8wUbz7H3DB2hJftScCUeAdswBsfAwOQNyoGTv5zOPxjwPIwo7PMfTRePdVnFJ
S9exvf1XciaPOVXMoOKm4w2wvwrDu1cMc7SWjxYxB9y0RGhK2mRLToWkkP4eZxyx
/riHXtWVYkRuwUY6lqra//FHZ23t3jQ0JNE6dBJgrLVVI8P7W8eUY6T6/l11JKpi
QTglnAcMM5uOCsJnDQ/etKe2THA83Y3Uvvs7cnS7tL8s3uaPsd9oj53I6/b1hiIL
xWec2/lnt9pWMHkY/jUIjI/dgVv6qMzuJmd1ogaIv/V+0o/4hgQfzFg7zni3hX2y
KmP2F3NFNMU4EfhTe6Mrp0lsAZWWw6VUeQipu3SIb2cJkPurQUyYgh5zmFT3av8B
WZ86HgbvlHFzQaiQYIX/bwWh/4odZaSDgHsmo279DKGumTtYIEH+roTn4Z4zWKw7
XehR0tqARmS6CeaiHhsqv21YcxapOCM64k9XYanqkMVo8xJi5KBE2mTBVAHoI0Vh
X5xAUTJDX9i8HMgOK96A1LgB1gkDOSrAPpoHsYyYgCv/Ereoj98tHaP8TiBF2aJw
CHT7CTXvAOFiS7fyFO/GaVBuY6ysAy/r2PTAe9zj/qv4FoCo6XYHBHXwwTNJoks6
eqIvs+OjuvD+03dWss0IxsAe2lbdzM78giqfszqM+Ew4FSDqgIb9MPo976q+T7DQ
P3ofR/Hl2D7prxTvIyFXfo7c6k6+2rkU07e6JKccYTNVguOtXqUl2Gq/IgEtpINU
gCZbmfGIA4PLwWSfM4TQn+QVravT1j3dYT2+QwVTDL66pQ90JsFJhDJ92qrShPea
FX/667SllBttLDti1oI+8I30wDsTNxjhUvyIDSZ42SLfiFAhCLZGcnKxI4hzfQUY
Mmq+NF8RtgwOKIv69b1fL9H4lCykR0GDmqiyZYbMwdSHaiUY4qxdINfYxnUANZH3
vkNulqLh53+657nC9bj2j1eOCXikP+DPL7tMruW7SqfaIF3tdzFxLkTZ4xjdLnmm
jxTQSVHuOj+Wqt/pH8Sb6FP1zfpiSl6cFhqPIbDtfyAKk17IEn2vRB1Bv9Vqy+PA
Plo+D4ZhOHBelkUsfjlQ/59SRMpgPQWCpxY3wZ0qKhd+y6SQU7fqEMUliq60/Rdh
aeBvSBc8MtnNRBQuvz1UCnEuJwS9XUw4r783p8HAtdQhUlHTMrTGfMi2oxcnQtz3
y6udbVcDbuBhqNosN2JPnbmyEHTt1pge0sh+O9M0kxOHZNh//r6wYcIEqnhD7mj2
A5YmfAzG/NvTPfIo7o8uQX7GWU3U+1nnFnkfb01KbSPFBWKeNULzv8P6tYZsvmeA
6HcoqggemHhQNWdXiCTi1z5bkrRnjiQsnqVeSgZPqVAjjoklvHAIsujL6Ta/QsJz
049dcNvMOQjeg6GI5/H5GmFFg8TvjYocb5GK14/Uqd1Sg0JXgh9WRz1W0A7tLM4V
cgBqw6H/eoYRMwtYXWisxKVZEUyCQmwCtMdbjnuUWAdDZ0D5irap3JOVLs+oLbN6
u7S/ZUGsoGIF95V8noE7BCe5I357DaY4+tqXARtpOzbTFXPdEGg1avhM7fk+w7y+
EANP4JwYo0D6XFj0351xi+Gdtd7W/43XqcAj9blJy8DmNSSSj/H/UM+A1MD6wnwG
7Xf9+5bL6IlwtOeh7YD2EjTH6v7xIF8sj69naoHiOUy130ha+K+upIg6qMSSyK9t
tQSmh7cT2DXSCSF7HHkYo6yh+o+Aa39kaMByoIsqtbKoMAh/BiFtbvBVc03AMRcN
dY86Pbuj75F+HzVCyGM2YPy2Oi32SteYDZF93LI9MitWIxX7h7ZkV/WK4bdcQ1Dc
fLZ5mpSDzNE7XyCS/W/5GrW2om9/98tYkeZCuyUB4LNw6hSr6JcLo3yGHhPIL2H9
J+VZxFw5puPKTaXSDPNjFCss7j4Ol9wREwp2zcEkfkrNB7kIbNyFcE1T6ZaYM6X6
EnEVdMsltbGp6xgu6g9JHjWRLxs4Rw34B5JPvhelYX96Q8qWpcbz0t+KxpvqnoTN
a/N5YV1zIrNEHJPWtPHYBHZa/fhtgCEHBdWgYlMFOjmOtOMmSva2sC0+SbpC5jsV
X1lPie4I30s52JFQhvUMumCPKUdjpf8Bx77hCnXT5BX5vKyDJIAD+TgfMaiNv07l
128ZXiaIUK8zakOKCyA4imPPOPAPDGDKdnbyZGB/3+mKSPS4kOhcoNvY3Cv2plXp
kDFoZ3+NQLHkac5KwbDgJfN/6hoE4qzIytpD/cRBSEambZ2jqnoEI6hSJeIZmiQu
QfKTDVBdCeSzJGjZ6WVJ/+9aEEExsfwINUGRbvHp4ZNDbflILLtHXy4TETEBuO71
akGfA/kotjUDyvY7+7eayjtlakx3+66CsEcoGJ3Tn3J2Yv+pxdNegAUv9NvyrUnt
RF4gJgihty/jMLjTnOlx5iXgpR8ZBJJwM6CAfYE8MhZc8hFOC6dljVAitRWYzbAX
h733HpelDJuqXCmpBbzFncWxxIIDnbzV+/NlTmVZE+V04hYu/g4lx5cWz2DCeEFU
kqBmdACirLuKIKbPs+05zL33rFAtySvYoOudRDezq0lV1+IAtCSQeF0hqo/REAiJ
UvttzoptPJJ+uYoaOuHNnun+j4DUMhxZKz55agi4QIzR6sGZ7jVBcSOZH9v0SJ+W
LL/RCzFnkHba3WnMTH4qrs+ZwlDOyz8jnDUjvoBWNT4zE3fvt/D6DH0m8p9Ymrek

//pragma protect end_data_block
//pragma protect digest_block
18jhro3rckj9zOf2ybBs9qUmyas=
//pragma protect end_digest_block
//pragma protect end_protected
