// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
sxRFxhpUeyZJ4idtqVZ6QFICTvv/AV4V+QtgTTkIkoctmc0ShuJ92u4g8r6OCfWgdLuAjHPpeaFT
g6Q/0XbAYkgxPilCAs4MozacskIkl/OEvkw9fJADKAzbF9TaSWRihv13BacLzC+w/nm9l1nuAkxq
4MqBnh6G8PGf935ONFNkmgwZCFCUZdi8RL96GvOlhJ8l8P7Pg/uQS79WXP8oBya+URE0xp7YN4yI
AdT/qYBXMDbnynxdNNxQhAFDVvj3uOolGjCfi0QsdBYWnC0O+DjYWi/QDCwVswdKRVFZbQoE9f4N
edNbF6o9qWe+p7GXNzlVOTPREgtk2HHRu/n/uA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Q2UkYWVBmksDHUD7aaHICaw5QCqi/dc5zl4TSPVTuskuNhY92/ZaGIZbikW8U1kamqGeF7KDRX8B
hHrunTokIxkvDGzJCvAKY3FeKJpS/9tvVv5amul8le5+vEL2PGnN/GU9QFne5Kxk4m3YqqC04aEX
qbEfdPlQllpyPs6sVgKFr3wB+mE43uU+j+J9DUnkGdFfrNX/V/+lkFfXVVqtm8IZAVcnhHJ3qOrG
JfQnQdsQqC0SydKHRy6oeqHoHK9WRSXdA5MlU+dQnXH0zBvkTC7v2M1S1/Igwnm8t3sFV7d+/lCR
1vpPXSeZB5Ijnhxk0zHsrxWMnCizVmWYiLzF8veKS5iLO/BVWaCE9As5Th/I5yszVlN/63I5mwqr
AFg5gig7UKYm+nH51guww0gv73/+ycPR905mpkgLbC+YNngDtI0L4l9a7k5t1yoYa3pOpoq1TpFF
PGnkRCz3Sr1OF5FIBnpidfLMlxrTFTDh1QOvnbUnXIVC5hcFB3LNfY9se0iNBa4OQaOeBJoS5ivS
DlT79eYqJv7c9a38IO7Ne78fQP2HX3S9Xh1MrNhxjfWSQuh9JrhJOWmHYN5+qLhsapf8XpmAKR7n
fOj4tFZe7dEs2RlzVBMbk1NpnFYZbIhNL3Zm9utA0AYnz0couxV2r7RIouArC3hO+cRjgOxgKJIr
WO03G6r18U2P7OdfQ990V6u3h2H8sZ8XDsFfcdaXQ9q9XfH0gSahHC6yqrZPcUKLot91J1Y/nCj2
m3E5tCd6v8AM/gbXWoAAU1PkrAFff2QlvtDWqRS3HOKcFRVKswVl2A9DwYndZ1eEEkeIWohuqOLt
FGLYrgnAToK72yuiRV/+j7B6lnje/5bULCfKIP5LDj6PsNMnJUmoxaAVMphi9voFu7cZPSpM8rZL
y4JOCGzE91R3Z0LTgV3NmHwKyX6lL5TVm4NeWIRD0lIwvgqUXjqcL2PepBgHw5ubiPfPIUQVhPbL
4A8Q6PRTB2gKEhcVmbX6DEHTKL+5XsuanPdJz1Sup5zy0iImwYO/uG7+ejmmeyMYBAD0ym0AU8IQ
vTXb2M9K9XBH1q1MTSJtfInx5+YMcUpIGEzDaybwgxH0Ioh3sayIgdgBlkaiIHreq/jKm2K47Ie3
oti8j0uBC4pC9iA6iNOf1Y+WJqKq61Ny9TDj8Il0YVA4/ydj4lz5a4L5QMU7sG6Q4CFNSbd+UXOk
Arq75IfViGrF0yrZcd8qUkQDwJNCMZvfQ7l2ZmydN0Zp+ihFL5hFsRtef37sp0/WW+XL2P2rLPdk
OD36mvQhVsF09Liuw6dT4zB1pPsyfVOrx5mMfk5XDEsLZo8SJ6rdiELTpVt1nwMMEbFYkh3G1y8O
EkaEJGYAZAaCdlYLTn39T8VUyRREiySY3vcchdewiWAp7XO08yvwiUM6wc9hK/h3ccsTF4+krIyn
2/5kuQezZpC+UBRjH5TMWxbTEF6CkFiZK+BIVlkuV4bO4v3J65y2qsyYMCgsmtY5F/2yh9rAtitS
CD9hpb9Hzw7QqvatMp6C/2Ks3XXKpoBSAHacbYOahSi7hIlY2TgPCEC3aHmzQA8g/H24wP8i0ykE
hipJ6S7H+A3JSCsu6Vy9NaMPV/DKQr0OZNgHAI0hEgTyd7uuy1rPOm3nWWZH5nj25Xeop/08iO6a
ytzki7JAoj1XThGMHHYKeot4lssWmoYvbURjHiu5YtBiGCZ2K1EEaCm+9CoA0I69pOXi/sxjV1kE
qtCK9sVH/VbZjz+EaE9X6PdYcJ7uQ0UBSMRS+fAaY5e3j51XzfBfxhhlGJHZkKlcc5cv2dVJaOIN
zh0u1rrB3npjtVZnwx6r6wrJ+COzQiq7U4bJbK77HfTQpNCB1Wt4YEPfwM8eRUyR2wI1cAgbCNxX
koUGJeVaZQC800XAezjRR8XbBD33SBbqJAk4UTaZoMwJbEtjrc86DwZxozuoW0ls5gUc8s2vBso2
W7nSBrHdIIYllvJvgQsP9qNsX3uI55NfTvHCIDoSIO6TyQW3fJxQ/G4Xz+9hEpBH941hdnuC74wl
NycDGFGYIzamY1oYLr+8YC7KMNRR1h7joah8Fh5hOSravO/Z2M1UfbYk7Q0glINVFdFOmj49anD9
/j3KSFzDdV3/gm0jOKSv1/CgWn7qnppdQjCg9EZhOliO0EPc7i2qk6CyzgFiH2kwNZGfL3I3jSJe
0wxbvZydhK9/pOQP8JWmLBIz2z7vBpG1auovyrN1X5zt9b8UQLoUXJu6oaDknVF88RqhetTQq+V6
uWGNQWG9+CkOFxGvBU5JMDdCdtTaDjBBu2CfVfTXHs/LOlRLMNrVfyVPmbbfZO/IPYu9giQ0dUVY
o2LjEDWMzdq5MHOaIPEwkqUvsH8g5a1NolCkbdPrCIQHMhVac+0rA0UPP//Pck3Y9f8BzUpYYYTk
7RSclIOMAvDwHImIKxTyFv2I2nqC+XVMAAdPVKeHaO2wwZoC/qBAcULE+R5LZnx+9x0s7XSbxzDf
ZGZ/SbvLBeKZlnMKkHmm7mjOw2SnKhz4+90gx4x9mdy2lJwOrGU3ybnUWi4bQkulocr4FSUBVAks
FKxHVKjICKun+XgNz9pdmKGEHNRz89qMLwO34P3+IN3/eioHXkMxzwFKh7AKy4JMyvev4Xqdd392
+B5UlhaWOD4BgYo4as92H9IfRk91yPFd3CGrfNpBo+BrAHr6DFBaplDPPClVm8YDrcMjJUIl2HYs
AwvR1WGlelaSd8BEt/KwYsHYm5kGVSJZNc88eW0Ymv1Z2qDNFNvwt7ECp3Hshi571UvnW4NOseLP
lS9/XSFE8SVhPLMOCtdWZb50DgkWStTpPNOHzJxJ+m+f5UO1m7AUJr9GVHbW3LKkjMXoKP4rjiRs
s0DuyzvuEbXgQIU+NdqnrfHeQrYpuCLsZdBAaq9hBiUGCMk3xFeb69qA+bvF0+F5HvzCgnQ/2E1x
5JjxOJQBJf2vI1tCKVlCMdf54VjPU9NK1c1Gk2vIDFFlIPbsulA0rzAZ1w2OT9wgZ2DIeuZjkunz
KxYKCFgxwBOKcaMMdjw+DH5T8gkPsFb8xLaGNwCPa54phjA22bl+oyd67ThdVqHEdIt0fVvkQf4/
6T4k82rnGSOzorDpxAZZbpwmOVPCvAuvtb+4OSW1BFAikBpl9R+Cs0ApAOgo70Cmm84MR0eczN2p
m3KQ+Fgm84tDe835KfTJBOEjnsnX55EqmXlhO4fnG/xlB77umxoCBa6pUy4SLDJiT+pwZ2mZ3BC/
R6qWNop3AZQ770yE0r8Y/C39SG3BghfIx2eWufJvBsX7yZL7okFCuj7ZdeGeXIEhS7nhUFvBWGN0
kmnZymdcHu5ufGl/WvgAY1NdzLV8IbEfyg9ezmp/v6H80Zd5ab3scE+JaZVCEZ79cmhU6pTxv2m6
hnJnPKkvUyFQmzqceGCJbqikEH3ueeugSdaCxTpMY1H6CrR7X93Vard3qUXrg6riOWuPw1C7St1J
fL7ZmY8CTzE2Xe3I9jOO7AVWrmo8pSYYYyqodT9hjJFfsFER+jTXAoHqYtbngnpbjRbMJwVvzQYO
R7EqRqV++Pm7a4+ADCslAmW9oOkkIkDcX6xhKdi9Sm8TIo/EMZLBjU5Lrc12zjHYo6AvIBFUQLvm
gfcpg3bMCip2Xbgoc8oqNWirjGms6lxRRBci0G/NeGJot2UZO8dvJsOiq/qX3lW8FPV0rdxq1W2u
BKZu9gHzCVHwUU12ohdh0FpPsvlG/753cOi9aadXwuLZF2cxz3t9EZes6IWD39viphNgxQNYqUSQ
qME4j25Lbh5EzWDz9NzUYfJju3K6+5jtUytT0chf8ZwclPagrZXZuoWQYFBkfZbotQmG336l9AiG
SU86J7xjD4MUfZ1uNbB3zDwVJ84t3r9A+xA7LEGFgXFCwCEjfVRj4Bqj0bQoFnXHnx0Xepj7RbZa
G16YTYtAyap3f94mZgZMKhbJj+u4ek9A3xGiet2cXQznlr2DyS5q+mc1C+oBoOYSVeFEC9do9B3/
PaiTnTTCaI7pXpxLq6UxE1+EbQOr3dHq/AS3WcN8ddB3lP68GLlcWnYrvH/gELpQOtodAtDKPLUF
8YEbTO465yQDii9ock2pBA+yx3afiNLUy2jRovgBdusZKexvu0XuNLf30GDY1RM8n/2kCKikeK35
p/gTY1MCABXe72fKHBLCCb81s5xYtlrIhb2W9b93lo4oyfS9M1neX2N9y27AZEt0zBKIsBBa3dqn
7IrTBERv10TrYaVoYeW2AtLBmzaaApi3wve2WlMV1HmtFZR9UFCnST2uK2LKOqPG54xPzhhx1Q6j
g6a2uAIZqWs7g0YzwxLecAEddITfW5xjHNz9zG41f+qOmY0qXB1USqAG9vzIvl1Ukjaf0HAkwNsC
wpeLf9IyR4WOsMUrRrBegn9wowvHsz8ajT9OogXFBbTsN6CBhTYEpq48aL7lQusUdnB8BbSFhMoQ
q3yGTrpR423S1tqrYJNbHRVIpS0lrLbIBua2Zr8Qprw4+uSV3Z0lsGhbfRERrDkVYpTtZMzGcdtX
8Qad1SonFwk3AKQlKfotrNzFbyKNsnPXjNzI9qB+jvHCWwKt+4EFh/UIBd3DG/P1/afBwJrokk0h
kXtx1InUMR+FIV5/NkqWjZqKt7HiNXbQURf0qTRVQ6xNGiKYqEGMa6c6qWW3bor/NbLm/UwJNCAS
mV6gDiOuGYyEcpiWBSz0jbQzVz5Q1fLxGJXTrYsZMiA73nJffdpFH6TFgSgmyA/okACs363pXstj
9dZIK0eWz8/8xh16d0DdBCJLV4JVn7Ryl9tHy+kaVg2pQ/PG5LyqzhNflBQpl0g/A92Ws8dyCD8j
9a4kkytAr1Pv1ubQDMdSpYFmWQ9eRpnbq+66mxoz1UzckXFNs+tSoCFfXqzVmZgn0CXDXKAleL4Y
k51Rue9ZWLFwK0nMHK8itpCgPc7mxRQG/zXtqdJUUSvD30Kos/aOqyYcxUKt6/P4PtBaDB7Whb8H
WhNQKEmBHXwXvmYzcTfLxJO+C7bND8yR6YDo9C14Ux8rLPcAgWnVGKOHRKmbP4QxgUR3lF/e8A9t
ArZ+eU9HuIEwEO3ebBFgERT1T0r+Neen1zDrTBpkT3c99/SLK6cEpvFoXUpqPdZmChd0e8xFNuPE
IhgxiWgNRviT2CKjhgMdlYXXMzmJOP6XeZnU5pvZrEvtBKCOTsugZ+cuYznazceW4bsILQGsHMy0
sUpA2HmBjNYaMfIlfIBqnli+89l2G3H45Yc5XHhQ6q25vcvw+rkmJ0PQRUJlCzzEoNj7UnFdiyLs
JfMTLd2KL2ZjMQWihIRBWWk9gJ5gc77vGohPeFz8mc/9voNWgzsK26FeKWMmdELZnl2UCEnJ3AZV
YlOgpK+fm7T92oI0SqR0ax3pPwY6uq1wbHLKoltNlRB50UtHznR2dt1g3340QjmGk5fdd5RRrYq8
cXWdoC71yICbvPT3xSjtK4PB3oPFR9UQ+qy12BiBj7n0sD4jZqwjJhBzxGXw89BpOx60H5NZNweL
1/Q/i/Z3mY1QBbCGp3RLTSFyEW4aJa5eeG39xpNYZlc3l/80IIx857f5y9N4T3J0/V9xODutcE7F
MrQx4upEerchRK/cMFTBxdCELIcezqcSEBODeenk5WaYXVBKFoYbq9o5j0zPzNv8XByqghj090IK
t6gzjVBJlNq3BPGr+wAWpPrsltKdKd8J92XFdhiTwx89yPONrvdwAngZKBvuO9C+lnsIKCfu829w
RFQh8ifNU9nkqqKiepffwmxqOWR3kqrhILpWMCJceYaEx7FMDMZr+eKla7/zX2FRHgQKY7HAx8+b
aVqzK612sxVAuptcOdB2Drtis3gKcbHQTJHrfY1oaybq0jTeTPAyzMKOwvgDo24f/hTEWRY1RakJ
YdYI7V+eCCDCjbm1ixUZZKEvUyKUyvL02YQ4kxkMzeeFWzwYDM8rWQGHvv9hR/QHDUDqRd5ZHuOr
rxHZ6MtBlV/j4clwzPkWkWxNv+aUBUlRjUxSSe1vlaiKV4D2AipEceq26Mgi0ozEe25lYSQbJkta
+eI5W7Jv/3e2BicktO0iIR+m4UKIhxWmHwSHOoQiBJdYWXIKL6rV6FoOccKR49uZSf7fKDBPZLTi
WkYUajdgzkyyfXn+4688nhIgln6IO8vqQwPMz/IX3hGdLM3PkEFjDFhazP9j6cO8+6cN/v4lGjCX
jKEY4DMn9GIX7NcSnPuW54sktDcIAtVl81687c5jSw4fICVRTNY9ogx4zhzsa9ibf76hb4Q8Wc/m
Bs3wRwdfSBAsG413v3SkAfo6x6aPqvETLwZsf1b5hi7M3AJD90CQ0Kn6HwF18N95R6f4/G0r5FLT
O3k5GSo0cJXV9RzNZlcl7HBxFSsWrS5Lv48mA0M0EKMsBRHxQKW8juLU3xzYrMMq/fPSZv7KGv/Z
VipBPgbAIJbdI/HGXe/3U/V3/XC3H3T4Lb2YMHPL7/1JJxhia3gJJwcWWrDpf0eJjODl9XAoRcoT
ZopTsSS4/v0GVwqQARaSNel3Ngu9+TQJNGKCnN+T5Bubmq4TCQteueOint6ZEfhALoLzyV2h8Nkr
EnGVYRQivjYEmD+cRIxOuhFrOuasC18WiGY5EB5O9cUv8yiuH146FiVW9p4Gnxiom/42+2DwJVxY
xX9rOokCKePBozlY/oBxF+QQ4qNH0qxjSKY8yNiU7fdRLOhc6aXVOvW6Zkglt2Cal4CLnUQ6+vYo
is/4mZ6YLA4LjxwwcUp5afElIygypvEXPL8tSHDZTFgR/6xPSkuJRYw8hDTH6DSWh2lV8P2buXye
C6AJwUXGr/owXVUm4akBuX6dqeqmXa+1Sy8w/c7HHHrPYh0Kt5x0fwWoKswTjyd8lhz/OmEsEWYR
sj0h2lzRSiK7fU5+NkXC427JyqqkZoGUiyEoLjMLCp3QkKtCIcRmrH/ZRfxTZV6xk8uynJGq5oQo
q2m4KSOuWfz624anqTwwC7+RQFIP62EEF3eobrdkSJOTTn/MySIakjA3gMMCxIegPEGmFM5TjVw4
Zc5mFdVS4up0fPWXVfxKbKZQf+pR0IiNOH08l9A4JU+JGz4YHd25pwXjX5cr3J9dQi/9Tm1ZlqEe
UboQ6YBsaCVwLqPlvfSl485Yv3Ljm7qufvei0SdnrVJhy6lyfsDMYzw1+HYsYNtW/pikigjAJLNx
HjGynuU4zEdsGtRrhE2pSwrbSXdTVXrw2F5iiei5sIU92oUFom+sbngO12ovLnY2QNxmJ/nl8VJ2
2ilLxaNhwcjM6RanlF48Z7a3CE8JA+RCGLSXD8az3vDEwRrZvweHryE9ogGyo6fwS8P2ohKBh+gv
24PlkYFNmgVefsAvQCLra2nqlI/DGWKoWAAXwDp/G587ULTsgQbdc0RiOzLIP7fGZXLZXJ1QsfzX
vvVxPrSKJHnBMgTy0JOV+UonQDXIt3nKQoWJJTpZ2J+sdFALQAr6/h2nrUhi8e7Jnkp+aQi7qrWt
Ks/9Bvs9X1D9zvEbkV3GbSKkRZ9tJ8bam31dvG2dkhS+jAQ8+hYMJ+ZsLTJQD/5Bh+ul/HNV7xum
E70Dmsj+MRcR8J/bHo7WB3kD1bf1OaozEkjXUJJoScebxr/CR1KFzvrshMxBCQ2DtCt72ti0QBoj
iFEygmgc1itPZyTS3RsRL2qL4y0TSXgZRmVa6vhBv6UtYprbSavBlL+ybXFQTMLpvInogQiEgNe1
Dk42AEzhCFe7D37YM5yBpCLTl2ynvnnRrKB+qObykNfi1M53hO7SKg/I4H6D2yd0aOqVGKBe1gD5
ADLnjxm8m/jtfanHnkLNWaBaSBwbli2pa6+VH4VwYu4hfMD5KTWVXcsi1QK9RqEY/tKmTNtPytWw
+f95uZGMYS2w8TzD9BghJW5yZRdG5Z9UbuTJq9Mr7zyvK2a5o7CkDFjJj/7wRpDoI7f8K6g3SJfg
5IGRFURawcTZck8tgQ5O21S1A24T9BAONf/v0v5Zt/dnCyuc4pCFPYMsMqfERZA1MfaOs5Xb2hXn
f81R3azQxvkhM0+boe4mN0cbBDhjwKoqbm+Eu4r65LG/r+HpsTOc1VnLjCy/tUsFi2PCA+1r5I8w
WNItMNd5GQ7QoFOxNh4MIjCp3J2M7PsaCd6s2fCqmEv832ox/4lcBWjivlzgFBO1H1MT55SYt+jv
1jo9oYiVEMHu4BEEl5e3RYe+GnWqXYLsn7SLa35eC3IpR0RT16weOS3AbrmZyXmrj750VO8uFlsv
EbITx4jF2Ua6h9y/k3eAz5sQpyx5Du9ZL58XeoUH06ghILEshWqrpY8C4YlSUFOI5qAIPUfbadk6
mBt4pF3qKCzb8nNU8ETHTvct3E2iojysOiF6nPmGDOjbdAobRLEGUs4ofrN5qAWIsuBlnt76Q8aa
EpMsTivSp2EXFurVjUwUwsBqXOLi832sjeWGJE53DaPRlbPcXchfn3jOjz5ACdSV3xJQMkzEdca7
k4oQzpdQxRIWYtzsvQrJa8oPiYv0TzoVG3mvLLYYVdJTdtNHQSYDuQKiwvo7/36OnF48dazbOeag
vZ7SDiJAQVUi8Z3aV0wKNLKBfsHtRz4PQBBO1n6Z2qUYE9StFXuVnglseoPaGx6z9ovwNCmvM1VI
Gq2Q04y8Gxx6IcuDw9/ZzxcBoyjfqNzzOdJ7jW30SjzaRthzvhiDhylvIBX3rFcd6Vv+RC6kSrUT
NGvvoQB+SclZO+yrmWixuEM7qoVN11xv2dGbOz04buT9jpDPzI0elk35PJFI+0FjoZb2OsYiSfCO
XTDqBZK53V2/5/a1U4QlkRZVK7ensZ8vrtXgNO/Js/xI5/V3tWqwXfvUqtLrGhRNkF2QwvzobzBY
090F+XW9y396H0m3OSsp7SJAaUgfB1vTom6GBcxaS1inFoA3PxVDQ/h2iXOU7FbvCwNCUYfWAKOt
BOuOe2q7C8wXdBpLkqxMUIegmti23+iD+ly6rzZp9bn5fH4/pj8vALjpcGdL44YTD2AaDpPQNngd
f53fTezBI0fPAO6NW6PQ/QpoQT9U8UXxMlpEJDFLGc05hSJtzSaLwotKBXVPYs/xKByO8+pCNhKo
jdXloZtcBrNs1zmdH0TJlDfdD2KqnJSBUfnIqMSOnC23y7lKYgBUJxs77Sqa2qwkPZR6+PjEFAzI
cXeBBE6dY9CRrkhdnLlNCicJyRYVqaIIzbY/B9iCpbRhtHxPe1PF1umyWN74abMrwAxwyOUUxVz+
iSuTv97AwL3XK3gaA/z7R8H4OW3HRhD1QMdOdpwn6AOc9xYXKPZHlvQ10sVWcipuSkBctCFiivA+
7pWZ5KJj529psKqvM6+ZLVlMvIBTj1+Z4cdzdlnzGIDeSwI93yXoRprd4jP0/4yPf79nirAMTaKP
+v63GDS7dquhoDucnYkl3ojbD0+EfHHU5jt2FN78/23k4Cqm2D6mKsxSkYtZKXGD+TRo0W7TARdJ
+KN2et5tyecleO9T9lhEaejoRi0BpyfVysuesxu3UzHfA5n7zWYTR/f2ob698+2GpxRi1A8kG9fj
yzKG1QhVqwITcZVLHBd6ZyTUCZUsdpiOIgoAE6ldB93pyZh7gonJAKOPVZracgoS+60rc7rWuCJU
jAXon/lf8KJPEb966hurikd/r7BI/SxUiM7pjs7D7t4xQDdGkgFxr/lOAr3TquA540lsFv5plycp
7wWw+Wyp2dSjaIDPWw2k8H1qumdufj2VfCvSYMqmAZpjspIyXtccuqYzC/VLf4r+ezQneaWyOWLg
qg78r9SdN7tFavwpMrdiq8DpAIY14FgvRLsivjWBy9AQaiadThUB/FVLQIvPihE7mMbswQbghldo
3W63yqcJW+gwwzGhrROgwom28Gldlrh3f5/aNy3xfTj4Cg2/iKBSOJ+erLDFf9gUExzDaNwWgZ2n
Prw56NtBdP7lvhne2CQTkJK1X+lsCup0TKff211fZqUaidekhscMw7K7zwRmpuw++mL88p5yPC9w
Ie3aSqhiQE4LZ+yU2JonErWJ7v9EKIeL3hEyaCNAZNln5x+mEIRh7V+D4CAjoM6WgARYfZv2CDRM
mDAeCZfZNQrzhBr8DDWqaDxDAMbTzy5KsykG0cyy8/he7uzqSFFp8uWWUHX1codArOyLSZSaLEWS
C3hHauU1lcAfBGzy7iRTA9Jw2ePYG9ynhOH/ZKvefQFeo4BFyW33mE1gNYlFFPfxXHVJg0D44p5j
WUe7ZVbCAURQI731KwsGsA1iOGeeWUmdM8Yu3wYyNaCy4SJWH2eAUx5R7HzM0MeBnME1UJBrnS4a
QKuwrIHMEmnzdK5A7XRNjwV0bZHm7L1dWxkKOCf7fl59iT+S/uELq4TQ5wXQUW+aoO0Rbk5XSF6g
IYk/i+4GVyCljhaQI4n/RnDqvCUge4LCShyqdLABcpiw07JbreNgRw0GGj6EVxEP7TwBke2HqSJ5
N4iTXhMeIyr/d7BHZ4vqgX3YnZWC2i8P01scG2QXEAOJGciJOWnUjD0DLEy9K70h9HqgbftS3zHJ
ye2yD0Rpo9jeZsk11G89heRACtCPMg9qzDWj+8JPxu7+hMhquCBT/zXIG1RjVZPhUY+cQmFdOSkN
iEA6TMGcXFQ3YNG+iv03bQRSRcwMoL6Xm5DrS9vyb52RKHtMv+e1zv5rG6ZIsdct4FIS/onYozfw
nnZwya2aUjOf+8D7NeehmqLH79itA7U9UF4Q7uJUBkKvgtK2/qOGH8LFNhFC1CtQgRN2a1w2c0go
bdRA/eK+0QuSyI8sL+tP9UsVowQfYhD+G+cNZd5q8c5xhfoS4KOTgSkr5/987jY0KAr21hq7CnZR
l/6gVKM5Tjmu1xiCHxDGKTp3szDt4xxLB6j0xM6v7+QfQCgmu1F9O/+pJCn1Y36mfWIrwWyvvQI+
PWF8jQqzKhD1xlfhudeBtNcBVHl4gjkMjUjuhTIgYKvwTj+o1WgWX9bfn63js+xjfVpaNSV66mlm
+fjx7aPfwyHWJbBXPruHJaqodm6CO3+0CSkIKfhMN5xDyOFRohFprfkmxabY9SdQM7wL5PVK54XE
bYDbPGgjkCBJ4kW4O5mXU4GXUJgD6jV4aTfw/fcWsb7Z7/kQnuDdE/XAPSvRFlvrDgvDNWFYNaj5
no1hfKYaICCRisbpRIifqp0pjNGMd8t/9/dKjb0dCIZSarvMP/KgDqKs33hZioPVltYthIS1LD3R
PiB6knSKeh6F+zCYczMfsIQogfXYi8mGaW5ZSI9/wkYqe8GxC7WjuZeR+MLaEfPKMk04RPAdNkIM
H4C7G6aY3kfwFMYxaehL1lm56JdjYCI2NW+/Dg9v5vQUhbgPWJaQY1JkResIxAVyJtPDy4SuZHNi
nIBHAr9nJc57EhM+C/qCm1jKenqRx85+6DYZ9jfiq6/4TeybsLU0RfJ0T/2XYiF/Q9vR2yj4n61V
GbMkGnGNOwMa7pOnKAN0qsgywXAuL3fXM5OWFNDnRZoT7eCfYqgFEPPHbeUFDZEBkGSuALSfEB5s
2JissUkUPmJuxiSvhqRfAvvTZQytJHXpV1awB8JMjAv0xobJFVpQFvL2RcTfF+7xnHOXYsXGRPz7
Rvg3uT6lPehtidm0jhng0MAq1ZrDm/lfGBLAQLOvgC2P0FAY7gZanNo/OQa5HQRAfBGUCFlOMi/O
vqK0itnB3UOMU4EIY4HsHqrIQnlsx+58Y8VgLlmaj6Oma6HStNy+72fMKaU5KfWsjh/evTIVJFTF
J66cucoZW3C5lyMP9LIP5RvkIGgeZz79eIrA6XRB1qx8xQfi8rJZVST0l9C9cVClnuzqesjBnqJR
5FfrhFrkISkWJd5smV/BuSfH5YzhRicptNPIYSk2GoOXqA6ZKzY9JzK9BNaSVw9dW/yCpJIL3YAM
7vvD3lzgcms/kv/IkSt/SXL01P90AM2F3J3GlsxCCkCLugWa7RRkgbJCzM7PIZex5IspU29KaMvO
qvGTWTq3TTkxlgTkvn6aBe5OQFaJ3OolvUAJ9YMqT142Q+UHTYuaTwsef100AS7R3Kj01twFPY/6
/xUZ+C2LsC+abvL+4vQCcYLyisz/H+F0Zchc3ijMHvN5PQ4VVmChsDQnGeCwkh9kauVo+iqB8ECq
TJ8pjEqnGPbzbfAt1kiqr2TRp8VA1BFeR3UBB3XYbejVYEVcwh5KjWEl9fJr5RPDxiKVGC7WoGeq
06SmnBfd1nHDEdJxtY4mC6ljYYj0y9vqSAi4FIvs68lZu+ozx4Ds/VWm8JL56MBWIdOsFN+A96wK
aQGJEKIAwGwZSwasmkD4WRlcsSXMcRLt/bnZniZ0dkUoQNwuRFYPIrBUQDUPCvKb6eOXtLmKhF6n
pDuZ+pahLdhC+6fp0ZheTdi5kW06VInB4GjCQSTknEz6l4wV1qvBr6vsknZIOP+zrWjR2R9zgs1F
VX63awE9GdesyyxZ3Rbig8v7Rq2koQdR1wJg81uNHKq0tcx6v045CgnAD9LTUSQn5vKwZIN3+/wI
U++spbReJkba5kF+cl3CYxQPR75XBIP9sS/BDgcwp8BqsBr8fxmyKqP8A+FBHOkMOWmWAfYdGS7d
CdmtTiGRCe/+zffNUlQjDKtWt4sqcmBQw0LJ89Bi2Id3EKH0tFALn+UL7TKkVgVfKEG5RxOs+tgM
xp27zyWpK14itulKY3WwIulSZslTrGudlOhiGLgpwtAFxXvaRHgYXhvU9NihSjZhCqOOD41uMp8r
3njmUV+Voil4RTFv3qzglYnWQhJVNr794HB7qS4i2a80V58SbdmfVjFPBjkVDh1ppcWmpl+TZtYk
fv1qLHFChmlvntp71ETQ2WRh2b/iDY490JgBIPFQI+I+fwYoQQK0UUmzaEh5UK6+zi2xmq8B73a/
cWxq7++JE7qPwjF6nB2kjlO8yeZvKT/lCLOLBUVKYp0Pvfj9VLrDbfGKcrp5qNzceMHu3+SRmvU5
MGSTqs384KmjOp9+okLcLgA6SyoM1yZrKgzaOiayvnH0N7dgi6y1WKghp7H8hKeolxCBYY4CSiub
UeS7YlAmBlwE1b1KVm+92Anx4CkrjEAbBIs2Wtuf4dbNRN+ddYdaEfEa0DnN5oIPj7xv6ry+KnLs
Rhs7sFwllnyQmniSfH0S0rsJMX/rI54b3I127Cw1Ar3r/2+M9OjGJDyV/tGONMlxCmHqq6sPqmwF
fdBjx+4PbFj5q1iz3XeEehdcb5qJ7s7uBpi2Q0BFsjDpg+VMJCJpmqDgR+YYHoDr6aVHk3auWX0n
E2XSXmySO+NoAv1ThMIuTzuhhWx8zG1+Ph1HvboEU2gvZqxnMV3YAh4RPJVUW1Faz0nUMRJRvVKQ
TNVpqUCZCyoEAnZf5umTnojP1a43D2Z2rW8mSvirEh3vMQ0UNCIOBox8k8hh0+QA2yFjG9jSaGvt
YvTJnKC94DRrWCSvRqWzELX+cjQbDgBhJSD5YF5C82V6WFOSasRljeVugW+gxNwz3HQ5g7oIlfeS
ULcKt5WL1gcWpgZH24U1qpe8sK9NWjmqJw6DzjMekjMTA9eoLbg0ucRmMItsiAdzJpJ//LvpkeLD
/i8qkegsNJqPb98KT2y+AWmyKbeg6eKcdybxdhSPV749UqmUxLGY8dKW9vuzolJcKtR2oF2dxhVu
R7VkHgGMk6O9uJeME1TqNCwNfD38TFHPLi/FUehtRiIZmZ7F2pf3ywbcxVhsqYrYXeK3MbtCy+8+
TbOUzc+u+KMn6N3HGQElo8+ea7egYq36mKMqy9vbxspFgue2t4h3w0sBOeTtT/UYMl2GH7iCGZsj
ric9RrQsfDtap4/YFBi59VZlV3YLgcnuqMTBR1MQN5DsA+K186k3ZnLWkLeZ+drfQ7SrKKn2fB6V
WmVwsV0KET94zZVXJfnyw5XvNxwgL40HO+4W3Gax671IX1FdPM+AOZ13Zzsv40Y/OZK2EQ07aPvv
/kszvUcliG5plTciUJ6lraHQZM822voB/2JL5nwaGepeJJgX6dXkqXQ5U1kvwQ9WlM13dde6ye99
sOm6hhAujQheUxBPLlPi8Cjff+8j4NAPtJ+6+4e17YCJQxh8fxDYRRM/mgg3LmPuadHTMh4CCjL2
RcVNpLgMZpvLdkHCPssJV4KIZ9JgiJ8tGRZTpWmzs5DsWc77H9SIRw41nQBDMk3F2DwG5Dtqe8ry
iscBa9z8xr1uAndWkmdE/1nj3ESkOwzdz6KD6AbxFNsikvcDw1OAkiZtERiU9EoSfbqekX1ejcGD
ROBwd5Xv30TAlEfO29raSs3Dmclp9tmDRYmdzvc/LOp2sYyWS+2Fp7Y7JBeLJQIp5pDlD9fI8bem
zBZCvZZ1V5UxFC10C12gndd3JwFDySDxKn4AoefjgYpXaLT/YDW9stATkMps0Z7wJSN+HznoL56X
yLZz9tCNziIzJKDRmyyUhEFtkadNC1bHN0C8qCNq9PEhHCwcz+v54R8/JFgcyPgZaxxFGnLRuRTF
W08IKb16dxUxGFYyac7oT3hONfyzDtKdpOTVFOPLYA/7s0Vrxd7Jg2NxPeYxrz8VJyfclOJYE9iF
Z7u/9Ljc1Iad6348iZW30wkQ1m+Jboig8r+g2xtB5gFLWFQwdaMAQku3DbpkYQSl9PW9EWFikOEW
L+41/EclIbNgTu9WTWFHKfXOmC6PiOiTHoNMMf7sLXflUnfcrowGj1DYWZKUa2AdHqvivMHlZitl
5reKnHr4wPKR2UHx+h0fetFMiHadWY9bKl/odpArfeCtDK1nur4KjKIx43K7piGG0OO/hJP46VdX
+jdEDodaUf7/rJ5EXSG5xSR4f//bUZgfsj+KJjgQQoeRTsP5fXUb4onNTmL9utkCzMoorS8hpmoJ
GTBE7UfXh3IK5KPFffrbLwW4bbcitp7BLlxsaJgZ/D3k3XQ5rAJjMJ+oTHEn7rPetfgdiOFHE/26
/V/TQBVUXErwexjWl5HL5FA9zsO19kURm4Zh8NDyykP8GCucyw/DPaQuLZlJqVBIzL1d3ZM8t8Os
dUk2B2SKOVxRZl9TUDS8ZDljpBFAiXNVIkTSv9mxsl7kUqhFVahT4wQM+n+wDvkx0O7/E4nYhv8+
JCzGK5cMnZot0+pWO8Oj2klU0O9ndJHBz/raUPE1Azkr6Yzj6AnQ9O9EFOeHNK1T4BHPionrlkPZ
njmdaU3Yg+H646p9QWyy2vep30bqWQxxDOHyxUaXAUgqFc6wHUmo+AzXEYgD/xD91+Z3FamNRA9/
XjeG5YMuw2yE5CV0TabCARUGuxIXTATKQZBBj7l9djNdAvoVZ4rgmQQOWokQPTTC3FzUYDiD2sab
QFRBS+0mPxj6daAsBnWrKRH8ztXRqZV6jQI64D1sNoCht34deO5o71isIWx1fLP2jbaORkFouRdg
CaOz727v0r0WIFhIQjg2i6y4dRsF8hhChNVTNzZYDgofPotJRTEfHyHntVzxu3GYzvBwIbGnOmzL
rmdzIAYolLKE21U8b5+h+xiHDWIQAFsekObg0L49KYa69rJIpBqVE/O1l7WLnzZ33yYV6gF6HCmT
4WzH9O/if8OpZXkcgg1Ovh/v9J5H6GXCb0Vr6j1UlGYxY59WzkiYA+jQD8Wfh/6C8rE34GeNAy1W
o1fXim4NO76JiPFD2uweQvMrdNAB8HyEIVQ/oRoXdZSxAyz8U3boFE/9AT11IniVw+k8bXjI3bV+
shvgPsIbhzCiSX3itLag1DVC3zoWGArnvPlDCDSBmZJb5u32Lobfn+KMPhZhldF5YMwpolQv8CCJ
gVbJOy0+LqyYOkhW+Pw45cndMc8LY5WJL/Lj8V3lrrGZogatytMajGwFm64NCaAHHDld9Sr85t1V
mzYrhN6LwWqk5dBgOiaxNlagMmJENLBaUbFvOr0CqM6kdXSIDAJQVAF1ZWThNERq1gru7fU475Ei
AurFTtSYGsmLUxVa1SnJVDqAZI0qJ59afa0gs9asWX/fCzSlB0kWoE34OEzOmWnpYUP7OtPNONR2
He25Ime/0Sw7EJ4xYc2u6QS2vyIm/dq+Nn5ebR0MWzalNdCtbb2mha92AYJroNS/JfK6WszWLZMV
NYJDJc+kSFVU3ZvP75O2DL6KL6LtuoOill0oTHGs/RUtKbl3hjRgPC2dHUbYBDBPDN4EsTkMDPAZ
gfwB
`pragma protect end_protected
