// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Rb5XB5hRWPTzm4DEfZpdRSndVbQxUPqAAKkX9zSOrMlA2y3fhc9BEVAVL0qv/9Yk
QG9y3uhJqadl1VpgR8hSFN2Fo/5FHUKGt0NbNQh3iVkBqmnXiPuz+v6lfYY/GNMQ
L7HFD3LLe3bH7YYFDqzFhIt55Cp3QKFtUKO4NUWwhx/MUt2XcSk1MQ==
//pragma protect end_key_block
//pragma protect digest_block
7aTX//wRVyeo2NLSNFUTINrneEE=
//pragma protect end_digest_block
//pragma protect data_block
ic3mZ+rwG+lDWckMR5UNdY5lQLAf4/hCXBbBgGhFWuJGlc296PElC/dlcE6vWI9h
9yAcTrpTxOoOw6uWDUlwpknbYkIt+U12Bfx50DoICqu3EYAqLdkj4dK0rXEqjXEg
6Mp72hkKjLO4w1rnx70gg966714nunY8XSzRcDT6tb2xbkWqEbVGBOn+/JZRIn9h
1Wx7UjsdMI37pqHHvPPnGA3dm8LEdAhM4zEnMsAS+FG/wxmEoQNsxIHTDflvc1nw
1n3zYHVlE+ZdmJVKHR6dnWIRR1580qbMNLsoPDY9oVqNjXrN2LODpQnCSGkvcP9L
W+K/t+Y65ZborxtUxlqWWkCY7AzJ58Ln32teq6IYiMScG8pcvZi0MyXitUeRJm75
uYkY4Jk87XNIMroRsrSWD3aJkrXmSP4nPNV3OYbkaIhb1hX+EEuIT7Il54PYMbYZ
3/2pEqR2svOKGItuZZHARks9GG+06y20HcOL8wd391ZWQHM0GWg2J3t2cCkNJAwy
n3u+oX66N8shaLgiTY3SIbN4RM4c3g071rKAIsbWlraLyWXbEZSelznxNOkhfw99
kdUS6uIfo9/nefSvB+CsKy7BUgJDlhHagSbsAZ3CATeORIDfT2YcBhrMAl26kRU6
aTLJuOyk1RVsWMbUAXWVD3imNgmpfKRaZM2B0HfDzhBr3UYzEhEaCpQsSU6s7Bu3
UvUXbsHua58/QppdcKJOFWTk91/30JeCHHCgz/4etJcDsbN7pHspKB+Lf9k4pWGs
MU7iWS38w1K2aOmX10SgSl3s3EXACGj3h9kXFpVAxwybs4cSGBcGh1sjy8aoR0BB
gLZRqXmeJpZ8YTd2tS5oS4pubtWOpArmvTPAr5WhLmdRxz+45I4Hm5ixMmDy3V51
fH6GibprNXsS8NJFr4FclSsns7/xIQRgs9aN5wQHGfNiFnRkdWuQLIvDTO403Hdq
d32S5sDKV21qkIh/0tIuROklAnlbiepF1FdB1NDsIq132bLe9Am0+lceP8rZzi1b
DOrlN+pFA50QgLGi19aVhMRjj0M65JxWUBoP4E9V2X8EB7HUcz97xztOV22ZwU/3
6N2H2xPMbgOcsfb9YOttnE5ypKubiZTLKp2+u1o2pQHl3FO+ZeW0Htsf7IxI3g2x
Z8vWK1OmDAiF1Lg8rIML3hG17EQ1/p0m/nAxLh/ErwM3LirRmYjP5zXzBlrazBPC
KDIVS9fjUuBFK+OMUecCvzn72U/FQhtVTFVFcPCruWSbjuRu8YMQhVKD3nLhxrR7
sOp2Ganh1ysun0iMkPkOfYQtp0WRegDm9txUVLTwaQe1lj3cig+Ruqocwhp6aInF
xnDGtrPKirrFHcYNS6nui9AL3euHft33uK3xK7hDAyd+YKVVFX3PzpxON6i11HtA
FI9vWWYtY2LcNJqjQ41q90oA36i6eGkNXqko3nxjjsMVKIDaMPXhimUhoxOzfItk
mlO07UfAbigt1OYsMmL/UQk7+KL/EBIvn2m+ET/Z6IFGp/80vbgBA2K9arxnh7vH
Y2A+q0KgB9j/CXAjyBR3wqgwbXfXV0pHos9Oll6dqG6RF4RpB4BFmOBcdCORAVk7
ipw3pRQsrVkxAF5Cuv8ZGzkFMAJBS1nUM2QFY+QqWETC/opTwyAaQwAgFqPrWGmH
9gX3gmfioQwOjAjLmaeoZ/rGaq9vZjNubNSecrQpd+axAZVQpCvsHYwQyfg3LmzV
+PW3GhYT46Vsfqr5oYnNxihe42vHkBkspU0+QwH7WJqmLTigr4U357jnvgbWVger
ox2tmt6DwaGp3p+0GHLKivvwda/1pdj5qajgLig++vnKqEks4o8jFA56QKHk68u4
Ic6vsbOKif7IMT940rt/7U2DpRVsfaCR/tK7tId/olmUHZ/koJNEykQ6EPeNC9ux
am4uDf+U4TP8EH3lbfD+9TNMJmUgJi8P4aMOU4+aKW7/0vHfMwu8isGK6LF26Gzg
3W3zBOhxmNETuPYSvkziw9yAAVMgEB/i4OXYdGsYUCQGeVf7LJYFHwaLLKmSYQtb
TYi0IxauLoX6aN6vMggRAkmzD2GdetOXAPjRHbYAQCXC+67sNnmVt2w5WDI/NMPU
M1KMFjeTQ5aD8e1sgDJ0nP6fA8JiGU9Om/975JIgttOyUFIoS3OctwZAp7FjiVGx
9I9PQIhC8PTPSo70tgrqb8oVlw2WrQfnT4fiIl20+NFmYzvL/MmZxHryi+3FhB1s
AHU7xnXHYMOge/JDZ7P2TEcfKliE/vl4Jc5oy4QZvboDhiT1Dh0a31w34QcGarfD
1MGZfrMktXMHsB1FX/WlyDtIQkN5+H1NpKUQQfusR8gGRL9Y2YFbxt+u4flOkQV0
2bdUtJ3323SPkKKmWsHpGugT27nzQdelojpM9iePWhQh8cOkvqiWne6Zybw6ixbJ
Rd5eCS3asC0wC/Ojs5CfoO0ja4lqzSVbdzCbq5UImoRcaqULgqQpLyOMJoy8i8nF
9oiBpQM0+VAE222yJK4qL0f6wDC6bxAN0jXXBLHupse4cXSr/Gx+fW6vYgFCIbQk
R0/2WCepnJj2jcT+8c3NJVo5hHQDzJy2bJFgXpJGlGZjeqp+NHVPZGlLaQLyfIDC
KvC9R+uZ5ttvzfZBEyNS7TkZNXyY/2upwpDblfiQ4I/sfDxdiTnXJWk5m512cU2a
3lre+cQYPWgTrCGsfp6Zf5tJhuqFzBFViuBh878Wmq6+DWAp4T8EF8tbAxCdfQfj
07KhyOl+xXzNR6z9u3usJHTAApBsMEtNqkjebGyl8t8FaWPtGtm8lTDnHDafDbjv
1xiiK1CrMU9D2wFInpWzZHCs6LT5DfSwHwQfqjLvkcAWYdh8ZYIbIrOi3hH1qJe7
9XtT8ISiLHTg7N/6NEFGQJA6vpFTya8ltIXuygq26ltYqDJ3lDtudwl3DHHt4QMz
HUqzAnToiANIo1O/Ir0AfxoebQBT8xWvRii1N6wXULcndJju1hxnJF7MgSmOPmwB
Rozq6qbLAz8PdvF/GzJdw0y2zCFFzFx4x9TK9zxMopmaQ92+V4Qir415gYKP84/r
UpoAic1m2ZETSKcY75GQEVdWy38oXdw2UvSSd5DbRpm2FCRQJ08KS67N0bCYGbSZ
G0hwOxJ3jO70sWn2BNf7XtkIw4MJK9hC9FGEAiaq91IcKbJ02DTWHTit4ggpSKAK
VAx3xSMgfHBcC0dTSdoQE77ImDYgV2yEHp/GgQEZl8juzmkQI53quVQeZvZR7TZR
gisG6N4LSmjz9sa0Hl4Ks9z+I2j1AndIBWku0fDYDVaIbpBJ+OC54WT8qLFihl9C
P8jZVvrwskvXVjhhcOjoGeLiY/Et2m6xktVYXPnVAj5C7W1lYZOzGPJzkiKlhZb/
8ANQRXM05U+coGGaT2UZ9DLN5eUDTsLWz5sQ0sYJGoVGKLNuGmOPRpUh1s/s/hO4
fSNJavdR++dIznkjrVNMBKlh1YB98dvLVSZaFlcji6Y2b26GT960aFuH5GIcVhP8
aopnE5JupiJdNXqYL1mF7CBZVb47k4WahpHd408f1eF8GcdksaSULtgpWXnqph5c
5cl6Te1PNjkyuAR8gd3nQX+VWs/53t70gKCxCZK+tjEK1jxQxZwjdVMm3xV3iX8K
IwCa002aFP7PAzjCZCVGCuXhwQqv9JVFbCYc5TcTV3mlVJ8N7wO3InxdnNG4lQzz
Qw1CbmSPinr0Z0Zs5nwRklaESlWFQOfh3J8o4l9I49EIGlT4r92ZFOZ/5b/RiIu+
wRqgQeFGiEaEEDhyIgdpWdXg89ShtOLFO+1bZcFTfOUVHC+ChZC276VDxmGmS4h6
EGVb/Jrg3D42f9qNnlNraRwQ2KHCNHKiXr7T9tded5XBeetepcgGR7hZSqn36dx8
z88aTWXmKqh46S9F2hKngjiB2WO2HDQlSdJIdYzUCrc1rtiDgbq6mTu0ooEsKIPk
5fD0Ksda5WQSFN3Ap9C0o1Mfy7FDVN3tR5/Pf9c/yb8IgQN3P9ODpPP50TrHz5NY
3Js9Q7GvEAqeoZJimoSF3M+0sIleSNH8LbG/kxjAGPgBaIceBDox+i9RWYLudn4g
UkVVSNRvMGbtcN+w2uh091MzZxf4A6bqytbVrWg2wxDJK6zPhH+en4ns3pgt3lb4
c/94U8KhWGS0VzvmF3nupOqUlBq9g9otnUvGD7BrudtjOdtN8439drTeVUZYsnIK
7yjqyic+AcWYZ/eO4llR2bWH3KoIzkuEe9H++Rs9ZcgxFUfDNx/O040pLK+X1RR8
sY3H0smVZgFUQ2JyHM0nEpXDKygf49FjWsyw9XIoqvh9fcZeBT1KaAs0xFNBg7Fe
/fANue3dRtedFCpXspmiAzRVdko1id1tIKxbZNRkF7+WgQ+j4GPnjda9FjC2bkwx
2xjacPnkrhmY8LmORIpdsna7WCg3Xz9YuTXMoa8t82Lv49awYSb8PGRlDF/Wnxc7
Tnntmx8NK3I5Mt3aa+Ewqull2KiLNCrdyOkROlwMzVOebpTRQMyG60gHm1ApgQXZ
iCq0sD31b/BJHsmFuJbv28seFlaCknnd8K3f7+9zR8FBTyP85oIJteTOtrrrAX5e
A6xH3tbK44TScsWc74mqfyX9wNUPE6/JJhO4amHHv8QnyxAiBm59GUg00mXLJLHX
hUfVjIQwgG3H2jdePXsG80OPFY/Q1LgVBMsWnulEpJwmO9DaBzHS+W7DBapbS7Ps
qHgGiYaQcf4YA+S86o1r5riISzvnJoFkcuyoZgzKpCRHh+K988QcJK5pe9I8u5VV
vXUdN7wd4PfG7MNM77OYgxBLRWYclHOkyb5pDH9lJWshw57eQylgmv3Duzp7z76f
u+DqsjB8wzjwqx9ZiqykHEw5UyypUbygM2o/o7XCGyDO2PM8RBAoEABUOglbtHtv
+p5gjxulwlpb36Qxwxzl7Ejg2+r0lMhWVbY7Nfd95KRmgx/K+rIiaVTcIGeX5EVM
G517WTMX0LP8h/ptCLbsMy9GJOAt6CChtPQxV0Kh96kJsa8P0QhGZFKxAip4MvE9
sFit/BrvydA+1FEOUK6ShXBNG8/sazekCHhCUcqFvpYlBo30ZSBlVY/K/jvQOoVG
ykOKTSTRRZqgeoVUMuEcomek02FSBW+UJwruZb4T/8Fjqm8Hjoq8RsltonFFp/D9
IkVK4l8u41DLG4yRscdTY2twj2D0bkKcXbTavtutHgCICRbc4X5lqTyXp8atAPpI
81tzthA1RYUb4KaLDUrByOFdG1l4NBtnbDi6zkQvagaAquWppoZmi5XwnN2IZPHb
FgPul7OKrQxvlyWApwpFncwgvMzhDlvXWVrGU9VU0+JDxLvtUHpz1ocO20expIzM
yqjzdYt7PwVZM2618DGWWI9tBX32xP4BhO0qPcFOZNipoopZBY/esuULDRC2qXDe
hfqCj2lSuDArMXSzR0gFxRU9erIAmDh80rb2dATA5kptKQUSVdqUjej//7DvCnWu
UaYIyECjPgcmawu5D0hqSRuoV0z9zMDz/570oT5i7xgOfE7W9n8FGftBfiIGccsC
KQucTjbkE3pjOV0/x8so8JMzEyvy8IL5GZp/kdae9Ewo830Rs5axxzBMGBYFu4FX
wVEkRW3NFaoClluzYKhse8IVB8b4PeSiwHoxJqGZKpDpVvXrW+ChlHzfoj5LrEe4
pzVI9pnRgWWu+lZn4ieza1vECWzfuEECsaeGQqdoZ5MRhoUiS2lIstWPxwPCO/Ws
Lz40mfU216O9g1cfPsRUE6tV6p1swadJ0yuVDq2pfZ6aXMumOwcXEJe7ABlYiDEf
CQT9AX4Ns6QkaZUbKQlTN/NiyTS5JZeeRGzzfK5DrQbm0J/GOF5jL33xLw/BFX8g
/zWJtmP3jrZp1GOzx5ZlL2O6YBfXi7HGm2e7bDAPloEokhEopbJxu5Cd2bzV3iTn
dxhDlvxURQCDDYtz4DpYXfoejsCQk/0QxLLo2UCuQg/3QGp9rQAArnRP1GMXAv/T
4hf6aAK2T2wiSRROCVkFDamVbi/jaf0xKmReqppP0BejJeY+HHAVKGDmKYg3/eri
UDCt/W0Vey2dSA6zgjErqYS6xPP/xvaAc6TkBY6hOZtbrwZcaP+Ia1lzOvhhqyNh
5nTRgRzEigSz4HAwl4nC+vRIvEgVkBntlng5PrdR+7qJOYP6hTy8ANFnY7VTbqZ4
EQvTvdUUJt3wtGNCtD2k7d5HFH8uZF7EO802r9rrmhgnS53UGmEwrx+QHfRBJuHu
r0WeLvF40FnzWQO+DZwd8T47GF1ZPfCTdJvmBAZDzZtI4kCK+dU5cZdx7bgclwpe
r9OaDIZUUE6Vknh+v7usd2++kE/33+9askCaQs6Qc0RBtqYgd1I9qyd2tT0L2q5t
r70jM7od/bOIFlrm/b5B08w+lbeZ9pKY2hridY1mkE3+hnPGj73u5MDqUCN4z/58
bZFVBeEJHXQ5DemtAGL8v/omQ0BZyxg7kTPqW/CDxzv6oaEp3hsPcw9vf4cEn9YD
CjGjXzfEzWbW7hAN17G35Aj2QaX6oC8qeeWRRq4en1CBt7zEegeBV1loJWrlb0xx
dT4CNW/NuoUrsntpZkxOJo6N7lHd5mfg7BHP6AIcplTFOnSorNn5ZqiplQPGZZP2
W/JeqGgrIoA2o/6d9CEBVI9ft0rrb7JUY4wyWx/UlxouWpYieCIDx77nVX3Wita0
sxJz42s06YoB2tj7Z5iBuqxrpk++YRf69NuloMVuh2u/kzc2ZDEa97qUfj4wpR2+
XKhd3nut1++FHKZi1DDDw4Bh1Tj9lP0+qAMIxAcL0JQbydzcDNzCj47NtcMZpaCE
CHl6drYan/XZBqRuu502KBqbhOtUHiiXpSvXzDamIbNVBlc2RSOl62/g0eNQa+cv
fhAhuDUd4uq9Oo+/nm24bKXHx6q01ojmKazL7ZYHST3Nl3fnRZuxpyXOursWvcit
ufnbyiyqoHXDP0Y+18tg0DmXkiXuKx96VKKJiDyuJhDmoeTEqNoJx3sUi9udFMhi
s07lH/RO5R/gS5KTbmJRdmbJJHnLUEezNRbhebsX+Y3hMN5T+nL5C8HrtXPAsoUj
oVcew8gUE7kzJ5KgV7Mf7wM/t78Fl7DrtXPA2acblTHO5t5P0Iu2Wte3qcZZAilF
C6CSc+YTaZ0TeBDNSOxhR230e0mz2yS/3rSWjkwDDXlUDwBJkq6zckH0asokI9Kv
wJLwF0+FebReH2KBuc6saEhcbUSGbfyfy/qh2tIM2xepX8X8/b3WoY9uEIdHYuJ3
0rKQYehXN+/Vo1WYf+XcAQZ5DkaJo4cED7cJMAsEtYjEYfKjgoclCErdWZBEwvSv
4CaZHNhPp2W6yA/l2JlXOfAT4XuyDC3gi5Vh9YAJ8fGXlwslxHeYXXji3T/ykGL1
5k4ju/ZS2ycnslzzFXWCoWPllYlJoU1zn1tKmzGkHVDCw7lf7JlMKWcEPe9n69PC
8PICcxYIpENtfRbOgxrmwrlE3rNtkBmLlsBozat+ZBVEoyn+GeirlaNh4CB9KTuf
bxVt2BCmcK+4vwwLaAu6NuGFHYfOmNx/5bYTOoDmTshGK7qY5smYFOfB+T4E993s
+z4vaOp1hh/VgSsBX+tGoL1Rc+Y/8MU236/moWFKmGHuBbNt4t130Pzg8+Tv5E5F
8gmNvtPc192DPpHd88hr3cidM5KQy6AhDaidiJkImWSP6YsNeOTtIkNtf2+KjnKw
PrVrqyAJuX7qZXxKZMx6ac9TUuI+CuwNBJ5LyomOOMR/HkAbau204+bbfJfY7yXa
dMEyIveUQ13MKokLZ5a3UJuihGuKZ3hCf7Ua0AI2cz9Cg064gagMnPtbtywPO+y2
JKk1f3EnhzRy75S81e+Qg8YNeMIjulux6GSu6C7YhFWsK07cCfINOanE8KpDJrp+
/Cm71B0xq2xRyD1aPCADafRFOot2DWeaZlJu2TBHkWPiD7rZ00dSYv24I9KrrMch
95pwVtQh/poLzKeUO+bV/ET6biy+0Vk+GQ1Y69+izJkXqBbwFWy0Y07EV0wor4sr
DAYnLjd4mWoC5FRMBi+xOJg6oe77ljJfYQABlikbdwoBdvbo0oFU9TGIVzcGOWuq
PIf7L+xVQBwzlnf/7hViRXkakHotxP41oU3qUNvqE+wTjF4z6nUC42zDhaI7tdy2
hpaWAcUd5w9CvzHk6EzaoycsIfxMu/zSpBhCHoWMEcIezUKRwanX5Fu5gzh18ANw
qUNAHjj8m3F9BxORj2c/AkcezZt5RiTFGW3dZUlH+/8rzTm14brOSJgkVw/EOcdM
cDBhd8eR4vFDo0aenYJYCuHQvQnKpbTt5BjYLezDnaINvKJr0BdJLYFnhGE/eTPx
N8Ghwrwm5ZR3KN+T+aGmnt2WuC7TPwGd80DoR4qSIWA7Bio7SKmvL78KEyZs686n
um/0SXaH/Kn1RsmRtPYBkRj0sruEFKVdi5NeLVz59D+nnf44grOncD4CZ57qX4B0
8b9E72zQYzT/K1RO+bqDzfW15jJmLjKYUhz6fcp149s3h0bdmHtlhdOqPK6887pj
+mhw/Qu44a/8flGKQQbrqVkdKWQlo+jiZL/41Ppob6LRXZyOU5oTthbgK95H+zFc
SkywFdg9KWTjFSm3OZmBjJ6oH2qGpH7ouxJMSm+YOtrds1shoo6cWnoF7swuFIdm
gs/tzG6mQVHTB1e9HvoeLr2wpS5+RgrNfqcNE5Iu91wgxkcoN/N8oL47T65LcLwx
PBnJZIHtMJiWQUUR8SylOMTuET2JNC4cBW0UCfH3tEac3Gx/CCsGXo1Hz2AtTUar
eUDCTFsxlyTfuYgDGuRTeCFbX4u+vvkucgXZMc145+JIE37URcGNEQZJkoZdFF55
B5R9jYVQTjKPrSGcM/y1XHiShJ0DCB/piGHg36L0JCxnpm6vN6DraN/WJApjwyHB
xKQOZOQrySTj716Uahs8Xx/uuuMz5XFwECknQNR9+yYswO1koXQZWTnhBghgDFTx
QI+C4EejPw+VCQRC8aTt1Q/Yhz1sCy+DkgI6ZfgUbjBCAIsjl3iRzzYfYAjTYeTs
4sqa7DujUrzL2I4gP5aZQBZiRZO4TjhKJI4vNv/3OozsBXEu1Wc6BhW3eLllAEIR
WOKe7fEeEO7icGmILcM+W0ooqy+TIiqP9p8jExk9CIUC/vOZ8XS861xI8v1mymfb
hYePIPKfJo1q57CI7U7yVeFPCjM706dewqDN0HR0/VAuaWVPRj9/i7o3JMXrhqjW
nNOoAw8DU3mYOLy0phz3qMtXyCgJiKYma0EG+YwNDefeIUFBjrNWLcngHTrQu0iu
IgkT8XTscKCT3rzEMNFIQq6JhocivLLyEvJWSSFyUzY0jt0AT0r/9vON2fiHJJ8T
d9sI/WpABVoNjalEDDq/goekZ5mzwGD6uiUP8VmBBzOysT+9p5UVo44yLqfUpmSl
hsOQ81abnr1WclWOoP+nDptmyBFNKg1o46bqJ9A6+6Tku3MZVjxo5ru1mfc6cZ8/
JzFo7oDv8NuEmChNjUnWPvKeha6blICVMHbRKFcRW81t50sWDKHznlPVjCrTodP2
TAVVy+03HKyg3e/mW8IMh45tGwtpgnpsQnlLkOKlcf1cr9URL2Gg3wqvNT5Eu17V
vhk142JyNOFfvOj5wnl8laAbaYnHDdNk0mAyu6dFKxVsCX0mJlGwRXlTbOgbiOuY
Om8bKuOpDpX2R0vZewAiKWicv+t9NhUvkWASACyz6ge/ZtpcZNjlEk2ujt856XTD
OcT1xDpfKJzQe12jHR78PxHVMf4t+zlN2MzwjyYdrPbtA90kQD5jwrNz7GpYH8hh
fyYfUC5MvctljaY2rj3j/16zpAW/3VKbp5mHpWBPVj6m39oH3nfnPPYI7VOWhcyS
dAsPHWnFHKiAsB1612WOJdb+Gq0Y8t2aHqsa8AtacS8bQaYWj9c9KHQ9F9yOPc1g
nyQ1iLBpbwibhHy/VDD4L2PAbqKkU/EQ4hqFDMXRaVRlVZSQ2Hf8HwOnbevN4MOB
h19pt5TxPAufRPjxtT+IPcsyxlv9Z3jRky9H+kK6yx2rKHyQHIbGz4iXFlD216lt
8Cyimr09Dq50fv2/lTmmvWnzNqER734eX3giKzKbcH1jhM79ZzLWpwOFTYZ1LVOW
+S5xMGkaiVXTmGopRVkrozY/zS31at2KS00YahhZGK01SFfdTrM/Zu7SB5poQEKn
qfOJqBhS6N03QiC2GvuJ/jAs+DsKck/dceKxFjBWbJmgHd1m4wL1QsiMDfE8v9D3
jUlTMaddOpo+xwyk97Hnjnon+I5TMynqXqdciTOKoPdQkAnf2+Vk+6kkP3sPaaa7
HOjFmBYPp72bOhsUwHeF8aZMxbN5tVaNck2eCPiLVKH9Oz+L93GHG84J+srfgqxM
EeWNJHGtvmkeog/CblqiXs8u6dEixPBdazDtxYYd5Eu292qGFVd0TNCpEun1OSSk
HuVaYvnMuNrzyXJkqqufbFP/RKRxNABpIBY8u1O+pZhJdjyzWcGv58m1VI/Tf99C
oyDEvFvihs3ivVT18/IeJ7A7KVaQCjevIo8KA2QOfkbc9FtxORprX8Nj4CKxWn/W
bsiuoCmZsLK18JJZOM9A7TyktAa7mGhwC8Sd2nz2mNkF+mOTdBJ60QXcUpvDwYhP
7wAV1TS8yQgAt+C9FmkXSjxWbd+501S0M+bZMoywHNUamhmOCvB6BXXoOKMdLXf4
6gHbOuID06bBO3rc9x8A+qmZfL5dXUuJyVfcKaT+ydS1sY6dXTDsh+wNSrWIWdqt
1qieoRtQ9KoGZuGvgqPSWhvg7UxlL4Dxt3oSiMk0m//mRj5PwKZMgxQpI+9UlCRz
Y1LpTEH5OfC3Z7+aDH+VYmtgowFt6B8h+myOsXoFjq7/7dzhCMq9ciNQXVVp6BLX
5TIK9iVRXFgszGy62Y7zQfAkXtk1CPFbtoOjVoCZ06FSBy8crP16hDDqZhRJ/AN/
aMJpy1HjPejwHEDEThbDnSa/GKaW4tNddEdS4ntyDPPCa0KBADehwhG6fH65740V
8WkKGD1HihtOQ80m8nQ4mww3A7KH9A2DHq5zaBoTurshjp9d78gFYAhtXoBxnXdu
pKzyD8RibEi6XVmUrFavdEgs98zXxy1LLYfplU1NWXB/J2zFOFE+91GVw6pYwq0A
IoIpCDxaSXWcTPujN0GkOBmp+uO4yZ8+Wp709V2pz6YdIf6Zp45ipMF9M71fJNkP
nSPfkmDd402/4/UkNNre+FRIwKMa27Dw9IwRNt+klW8bpAcWXekOyf1VwWAjhdsC
mCGoD+uDzLG38LhFZg8LrE3jTxH5SyOGyQm/hVikxceeLHpJnQ3dcjm5mf7VzgwV
UfG/e4GCK4pkXXXT0w87R3n1SgDVx6gh5d0D2GxFAddGENIBuSE4RD2n+gMzDmfO
xuxgJhdfRh70UasU2NwbUjzmXwimnY+ncRBmMXMTuGHpt8dLOb4j7EBsTVJHGXQV
ktN3MMR3Q2gQlZ08b9FOxA9K05fGX8JGlLaTMzBrnG6N/VUx4xo6Tjjhd3YawXS7
Tcnjx+rhfZB+/Y7t3MLzXacg4iFmC9QVbt8AYx7l1WNJHdSAR476bjZd/YmYorKm
Weccmal9wc69gc0dAofMPRcjOuvNvXlJLeooE4mBbm1yeCZVP2V4yDNqNBieR/tL
28q7bEcXJLYtQQbISaWNpShodhYcxtfEumQyeyQ/O9Y+bEpVqxg6L3JnLkuyZzNC
ny+crRsThIzyLatubVqvLzV8R6lzbPfYXLtjmWtIiXct1A5DhIiMYyWb3zGCikKt
mt7cg6RrDMG9XsheONA4Lq5vo4+Xd+wVQhU4thBwxCCCzdgVAXxxiRoVxp1HwMZs
3Yt2GE4RYjj10ovkv8D9g0MBdMCfuC6ePhQ2AGRx62Ob4KM0cBfQtDw/hjXpnrRE
o8OenKEdC3AuM7V8kREgagk4TUTKkn58PlwyIlF34jzwpvLO38ofkn4qI0PU0COy
40h+YzMVcn7b14UMB+hIa6lkOlhQYnoT0MaEF8S/+utM8c0NUfT1RbH+KZR2inKl
3yBbQMcIh47dGlBFgRZfAWPrj/R+h7pF68Pr90PoWoOZ7434OjBEINDbvwkzO6fQ
f9bcSddrZEhq43+GSRsPap5G6+3VXtB9hUe6PQqlcskUKSqpoR8tmznGAnqkGxQw
CdpOh6HGqmmdjwpBU0ypk0TqmzfkXjUbSk/FFK1ylutBvAlUn+K8TyAH49QK3Auz
q7wnBk+dh532u7XA7EgEZhdCn2nIYhOHTDQeDTVJpQWrM/JGIqJQuEdGa42mQRY1
1w3mccLOxynwwNdeNL7ippQS+nG6LJml3HlKn0W3L6ms+JoiQnrd6/CV2gTHqQ1b
uKGw1/NZgO+LJCZSRVg+YmUfCKm2KuZ0A18S2Sh70IbR8DOViyg31UYPKo/YAdEu
KigqZF41LGQJkqXqfRlzkJ9/7qFJOyBk9YpOTBzRi7UIISrCiBvt6phQOLBTsxLP
CLAvJpxSFuaR4pxKK6TnLe16X55T9Li26F5T+F20MIp77wQhQ1iSWNOMHtoQTvmj
cy+fxhDZCnO/A15QZ6gjOFyDDhBFI8xS1YVsc2WEaUvWnxc0kQ9QT6EehfuKdonH
6uHw9CrCmx5NISpFmbRGssxkEg+Ex87IuwDDmx/opd7BrHFZrU77hCFoYDjy3lJF
dE7+inBlqgdpKZ1kLeDXK7DV6EdKz8VAOl8h9XvpHSs4m47pyLxF4E4EAU3vapIQ
myd0vXf33+VYNMHKotoxVg6KJteLFWFT3CojjdOLPNeoP00ZshLNU9rN5Q+10Oqr
V0yjO+dwRZ48wSqg7SNcb63zfgOsSA0ZJG6m5KA7dbDx6X8Gss4fGMYlNGedUDJr
QdoRR+MOwrFuZoqp3Hp3hmYQUu1z1YaJ0ikak6tbh0m6c8wgjxkqbbEs9zk5CwcH
owcTkUWUEmzUdWKqF+55nrpaxf+hjM87TA8w65XYO+4bG5T9MLz3y+DEpoDcFXHL
bv7KjzR0+DlCAOtJgVMHGZojyGXItttGYX77YwG4WoQkG7ghNpZKJleBdmzRAuBZ
i6W6G5jvQHLyIUy0OAOgCj/MhOecfCRw5IAnRatVsfjHONYnYgD8h1snaCPaOf6f
4gy2QVAqe9Ksdw0rse+U48PWqCnS9/sNAKYJOJtu3aTRfriYq8FYJ2BdJ/opKujj
WL7kJjwNgIAgzaQlh2D+Q1QeznQSeMNDCqn9/tANYp8EtMlTgT1i6DYAaVuc+CQI
pU/E5lgotItVCp8cuYwVLicvkHwP5P+ypn51RSX78Dkt8xLleQRxk06B3QLk91xR
GmAXSbahxJShEgGACxi+AMZvXZlGUraRTAxrqOngJsumRqxmgOcnC6GNQXoNgiCO
JW46VghUcH61ed9ROmGkz7DrUNV5eOnMcdfBX7WVFM80na5S8OOxmHQoQv2Dfbg/
Knq8cXt1PdKlmlqCcBpnKH3YVTBmljoSsObdk1ZEFiYddYXHhTS0G04yHZ9uXP4e
23WdeiqNfmtE0tQ1bZGE6KEZUH8GcWkfO/VKv4F7XIm+LwYw7zLYqLx0LV3Q0pzy
ym4qMCbTRYmGgPZDl3zwQMA8dLWVm8VvSGmn3YHtWB44fqCND0xXWJ2wavu8LhRh
kaGwjZhi/2WxelsNnEFfB00aQ8+p3Pp05zhewBi/x2lxHFsZkVYjph8YTX8SrlNY
UTaodl/WZjqHO3xlJCC/kKzCuW0LmzgNLzYryED60eQv0xeYsUXTRdGk8mRyWO5C
0WY4Cv/Mrs3s0VVhV+8KE4bcvyVNjWvDLmtJfwfuGVaNvySFyxbpz0JMAGjihw72
SVgxH0AGCwFXw1aiS4P35WoXt86eS0fklglzzlAyt02mE89deoOAIlOlcKUx4TBe
LXY9uYn/Nzxqqb7s3igUBVUQX6yy8ROfAgcuNM6h8LhqcK740WWz7WFfoYKx9rkf
RHNMPZIvY7c1m3l/x1eqAe6gZC2GkUcNy49q7dOZzc3SPdqvnAU+pvN/dSJx3LKf
w/EN6PJc+9xj3uviUESoqd4MZOyj+zDKl9Jzxqt0I/FRyAn0x5GyWsSBBUb559yR
43J1B34736zXVwJfqhm63Adp8G1SNzR8zTPbsjGZYefU1Mpesyso4mIjoVN3Asjn
Pwezs+69ye9cr96ArRb+gx5LoVyZCrXCeP7tJhw9PQznlsjaOh9qQfCltiJ+v74X
Z/HX+E+hbwXFo4vVA1ieaheKnTkLGQYOPkHbFcdkcKjBcMHe4jH86XmkU0eULLZy
SUjCsTAD4yd4fBZ05LBj6yhWgLK2duVx1jW2A+K++cykgjZKsK8iyhxNGfo7du9s
hJ2HTGNKiuCIC0F6THMvzrXZ3mUcieUCjkg2UfcSDI2Ed5kg9oXU+b6PE3kcGiNS
kcapXxUdd7vJIMCpTuVZOo912bJRuNSl5ccZDVdQ9iE6F0VqIEA7Z6NqBp3NQKPm
G634TeEtC/J1oU9xA0lNAvkeReJV61ntsDHvN3KeejMp4LRtUopnf347/s6ub68Z
1OXp9gXtApW5ep1TZ8AhwucTYBgq/RkIzkyeeUMVin5RviV03sjNGuTMu6kTan8O
U7KlCAYMU75z5Tbjsu76ZAdPK98GQsOS21emTx5ow7cHgYOeeEjKNmX3vtIJoIsP
WgJpp0lSdEkSli5MNkgUsl+7mzwzmBa1vxlazYUcTDtbevW8lYOpjck83XTp3CnG
KkI3J8m4L/L253w5Ko09g7zDdgH8094HC0kLFefJAwnLHAAKofb/kgtlDCv0Dywh
8Lrhe4YvoazgM1o8yIX2OBB7XRIdtskH47MkvR2fs9BMhqg7d2fqmq9vNMb/+r9b
dNyP49Zs1WFs0POvIUNAx7xkHM/xz+4oNAAy5TOIzZCCAEDnmIweCEjE/FCMi0q1
+mUdcxBXJrK6RiDM0rNt4WmQV/GjMPY6iEPmvYknnnAKyAaT/dgWTAvQQUrlmFLP
/ZouWdERA1C/sA1jBHErybT3ZZJA+ARpbVCJj3TAYhYlcSiXUTY0S2QMPeicerZK
IZUMe/oYIODyKdoSrl0ozmdCS/q5y1cql0W2kLqWmkIgyVVZ91aKS7EYds8O9YET
Bcrubh0baIxJryzDuD9nM6fdrhoz/18/AH2zvO8DLL7SGNPwDOtpe/hUkQYFf5vv
5rnlzO9dwrEXR0Uv4FASgQOoog/MDJskIFplgxUVln617VLdCeZkC9V+IWQQV07Y
gd3vUzibsXUhQctadSma9fpZrz9a1Lhv1qPPwshWL8mmHUr7aHctuy6JHMj+3Itd
CFSufqRVeahIUXEZsTKJDh9LkCUlBInKmOng3/knFkoakv0VLJLyIyCWI6ljA6TB
+2TJQfIISHPIIt1YjIWsqqVzpUgiFy9TTVgWdvxG5uB15U1PjEwg2IF6ZFn1kO7m
yB0OYOgyF9Gq7fK9DucPP3sw9lDjXYYfvH9VXPWsjjxLYtGpR7I6ayC3e+wHFcIL
V2tKhO2it6yVbUQnJ3fRm3cUtVvZzRf2FnNc1zY2g7nZgskFtQ6DCWMj36zwWtEH
pRK6cSHSPAjVJAYV4+0Q+BGHzHku7IhtY7JjIf/2DnBmCbBigKj8nP9ijdHDUPoe
pR0MiATgP4VApiGlpRmDyThNcohSqoCwqskXl4+io/LxOSeBnJm5VORYxleEY5V0
yUTuMOjTiykIQT6X6DDuuhfQVAxH/6IlsIrh7WE3D3FtCWFL3fFm+78OvfHITL3l
TmNrmz6Dm8D818hWr/hYrNh/lkvaYsbOMywi+upK7vKsTOmddjvvDBnQI0nrIwSd
MxR/KF0SrVyZVIwRstgRss0PYWtdTbtzWkMq07zJNpgeCFLoOpiAigR8rfgDniAN
Te7VIyqEOV0OP+HaLtTCFHirxTcnyZzUfeOgbBfywrUOVGsmE8GKxqlpVNEE4KXx
y3HBHABlcDhmua5eVX2ElmXtb3A95F8kj0OYtT/3/+vd4pOnJ2znEo5dnwzD4HMa
Bs7Eq3aviQ9xxcbHj2OyNZgCU/GYkbi0CacL7jPZ5R6EmX5lVbiV01Pl8aRP47nz
ldCX3tEAZJGacfItkpFo64IhKe+rVMThEfYSq4h8wb4xN08sH/LA+8tLBWhUqZpi
BQ6qPdGoRIzNPvFTw3qpmgSvutfnE/LAtof2DxZtxsTOx6/fSvLwjaFMcdW7mw6o
T3vaBm1HNiebvaN24EgrUa40SCcy7VQ+nI00/9iEWgqIhCaJOMp77wY2OUUY/IR3
6vN10WZh9FbjdzQ1STxAaZPz/AYwWhMe/F8pUKAUs3UswUZ/sSn8DdCZB+7iKWOR
ouzgWWcBIXylb+D+lW38zscaS8gEaIBekcbeP8UeizW8dZnLDB1o5gYjSVj0vtND
LkbFjMTuCh2dsvxypxtJME1HVrZOj6AyhvFsGMt04vlBVDFdIx7+MATeYnfdm3U/
Olfn2ig5e8b79O+/9dwqDApCtC3mTw7CEA50xSt9ywPoLPtmFBloTuenn+CzXtxn
Y04UzjKHlRJ/srSDWAUaA59Vd6km6pOaoLukjiSz5I5nDXfqducHXFOMt15i3Y1T
G/alFS7TJYz6c2TB5veLWYgwgLAjpdGT15PTVYIJQVyLd06ZZw9iFDaxqmGrOclM
GlDwtsu0XO/oPcVkQEpTP63hfFa5kH1Yy8dVV2hIK+q+WilK/ojOefScUVzb4c7v
bzBFLcAM8mDnNgh0Z3RfB/Yl1dx07joYeAOxR7JeDjfzEv8pAKpQQOR+EvYcPG0B
Hwvof74YKINqtpRxAJKo4IXIKxub6dEiTVxmkoetsUlcrPUv3gTgAoN95/rGRZ/R
IpHKClQ0IleUskAqTD7HkLl4c28IWZWjPDL6Dy3IOA8yn5PDmXuwG/Ka9r5/Llia
sydPcDAPrmmqleF7/z1xTwMlTy5fkGCK2PbLccVY8yCoq54tElTY6eFWzhFYltbv
Dd/Yj9qzk9AZ3COkjeq764mFwzIc1ZNJvGStcXuiB8x4YPNRjPSqMbyRqFC6UfOq
Nv1UBEGknPf3Aq/Sf9LKD+pdmsu5WqeKacxYkpUIFNNt6KwtRu+aihEoFKtRHlAQ
e/JK+UTeiXVziMuEdWlftwuCUXbi+ko0SBF198lgAxM940ZJpmqT75O33FA2HO+y
yePvvvdGWZIPXf0lXJFxdAUzbJukf1eZR1MAOK/Km56yhQ01TyHjMjilGO6xVW9k
CBL0MJPLL8DQeUSqKi8dDvL+Nb4+Wy8M7o6HoPN41uytx3Bk8JFTGVwGeFCPSaLk
SvhYMpBlYRMAjmMAsrlPWmwpKiy8WdT4h+ByH0OX2IIsnHHgHLxtQ3NS5AC9DK0y
2uBLC8fC2LuWy20c6wpqQ0rgufltT9Wkgj2R+cifW+s2arwIMBeCEocZuVbP4Prq
xhORHANkw4tB3wfg9/UDZWwe82rfz2lSR7q9n2hfFsdtZ/ZFy1RTNIeCDR0zWMcK
/fD5N/NpbWIf70b1YNKFn+Xogglru+0CZw2CR7aR1EnrWEsZ+qwahKHf7ztBLOLr
Ky5arV0iJXlYmJKEiVR5S6Xo1PqEKYRmJqv9QYs28pJ9vMKcVpXyNUqlQQIwe80g
LBCmu/DdsW/WzCUq8Yk9v538JTBHgnxMdax4nc1WY9w8n4NvorG/XcHtgUyYLhLP
aYl/yBxeVxph9x+wwROEELXvFgggQFl2h/oVkxb7pDuW7VV+XawqMYv2EPjLuJ45
GbvsynUTRDHWq9e16ZHWwiTEyLN+ymaHMiML4z56D9arIqcaEZg7oN23ddAUAkCK
mrWPXUKmW7EW7DolLZHAQzMSJeNi9aauw202/D+jlXSF/BON77tgpB4V5YJgwwCp
d5WqMdUf2BJh4lM36DrYp4Pqbh3TsqGG0MHqHLYRGNCazvwB3iTw9gq7Wu5Gc9iJ
g7sCYBFkxR9YnGLs73yr5xsLA2DLQBSi6N2868C3al9Cf7Dj+VEQcGP4JBihjnxR
MMuQu9BoR2cgefboH7Qe0J87craD2kUG7Z9oaCn2W0/XnEOAiKd8bVTqysESLTSi
Jet5nkFjk8XJXUmDOKN+egktZOKVWiWzatS7wcZ8vbO3tc95fYrqPNu/WjDdsXA3
1UTQtsiHYoOaxb8WsxlALCv7B/mpM1XIZB22qSi0kGf+ifuP0PhNpjYQzEywl67r
WkLNKZd4PG+2CflGsTyjMGqz3YPeddkIOchYlGjDa3esI8vJDFlfV+QWXNNAKGz7
KDIjNDjW3miiz5pjn9c5xi7J28BadCcSvZAaq01POD2+TVyCH3h+KmHCSjwQ6MB6
NJzP6eqMvoVpfb9zLw0nRpz2qPYF+gZmcHV5tEwrovDqiC01khfbHiRLg/G+SOPK
4Wx5pjGf78pBattAy46zQ3e1QhS21wuB51qB7a+EW8+PYw2KLWSZB095FqDA1658
MeCMFKy7csNGgy+3JPqsJlMnc/ko/9ExPWywv84tBC5nE0HfZeq9aF/hnqukvImR
OAK2T0rSzovCdWsNY7Nw/JpASmu1pzP5HHWzoC6ZXOuCnHaf/6FMZq6aD1B63HXj
r3WjH2/E+mfNc3sLqzg+IsWkPPsI21udrELoYXJjhTYMAAVAwlHmRxeCX5DNT9f8
iAHwcFXTX/apCODIdzKQWeNvLXqMg914BDCs+7X8ngXbAfmVH1hLcYszRNIf4yX0
kaPMm4Em3gd3CcsxbQsPONG5169ovVBFmBXGgwQuufD6//z3YnCJGRTkVAF/6jR8
321gQW6hvRz1hyOHc//XQJK2NbQ5PrOad7fK2boZLD6NGGxoa/1T+ZK32CTulV2f
NxcfpKBd0hOJeu5z5llGzj0GVJiWn367fgOb6FYhcahxX5wRhA+jAseQOONQsel6
+MYQFvl3to4uO4TEjJL2ajzkndoJI2oHZ8VY5MGlxisofoJ8eMkXu/xv+QkvfO2Z
YLKCgfs4DqboyZn34pBAS/3Z+yd2eH+MDXPpC6IS+3uYoRSRQLfEOJMUFOEORyQP
v8CNahkmFH6s3UE5DtlP+ysQHgNdDynRH88pRQu6bwLImc512/gyVfRNhaZzuj1F
OI+9LeDq4QMVu+PR9pWVE3drO6BGjPrcMCCZJA9wPYGfRsRlfyxxneazljI+n/qY
fxSBRPHhoxXjCcjrPAyUBMoredylmLG1gJ2RqihiPdoX+MMqNGGpk4HiBLCZVMmF
8EBuT549+amExC5DM3P8U6YzG5umHt4zHXAvsysRswv+Oonu92k7gZZkQbS+Uqh6
1IcDmR7aOFD74a+qGjh+q3ccuOJ0L/L0DLPmfB7Tj3K3vzqmFozLWHH3OyrgJryj
/86h7YOXGoiRhEh3X02RstLtLbpNu+dHuAxHRWF6GkOiK4CtmHeGZ3fus5iV4dby
4WhgeoKLs9YLPI1gLz5DKpoLsagQ97ndL7KWMmMAidHMXjeB09turpxduFvEvJQd
VWQElA56e0mQOrFnE8Akud+D4FH3gPJE3TETBLkxMlr66Re6cF9lg5ikvBpgjn8V
1g0bbKMQdi2QFvgqqretJ9Ke+A67RxyMaVzMkqXLOqIFpkHtTUt/5h8ckgoNaBgp
DjIKxxlzrWCEv5xpKlFkIhCedtMQ79i9dKRSMUwmriSM0Wz6l7SknpYufM/QOB86
vTppVJ2C1DvVo6iRRjaoODjgzPRsKE9Ko5JlGOvth9Z2hHrWKssDG2oLeKcZOuIi
P1NB3g6Q5D8G4ulmsM/fTLUnLZrYsramya9jwKFK4N8MgQmNuAoFItoOJsXtN+WG
wuXhmyOR8H93PMyQdDiEPK3D/6vjO6QtTfphutnOxyTiPz7MsmX56vpgdFLHpnls
yS3jyOlbaqGBdP3YjcrSKlFiwZc/NWeg/IimHkbdcOKQKX1A1OXW2hfoCUfjHgJ2
4RR7IEwkuQsc5HnjLQDp2IKiWYEflWBDrdUSeeCb3uMioOnjCeHwIiR0pEE6UBlM
c45vrlPC/XBFmPxtox1Sue5Ziw9IS5qSxQQxZkQjcODYTk1rJSqO8jfcaq/apIlZ
cr+h5HKxirjvInCeclto5lMosZ/6OhlU2u9AeINO6d6kFcBPSU2zPJ9lc7heJALF
l1uc8RtBZHvjmL1CRsOMfUNvvIxmvu3mNCBzaQvlJYJqIPbecWc46vgOMlmAGSsY
OrDGqQkdk7i24GAnk4PT/0w40BhWRO3PrQWnDya1sQf5Qt7WIcWKMeNnfp2za581
hwHU/Y/2dKaibwp6mYiQwqdJJS0UPLJORzgFJsLXST+gjIEhEi1WiUF6NEfa6auU
0UHFT5kze6LSI8wikkW1JPhD0YK9sbGwUs4pf8XV7LhIAmemrSGqAWYraaiQsDif
7xBcMfQnqemHi0QH0V9Bq4tF5lVLb+admUZYDU7wmP++XMyZmRSjlX5qSw1lIX5G
UHUW3rcDav6Gk7fKTHvJpffI/RD0G5VA//eG7XbXgQkRyOa6jrsYoBQkqaLauD/D
yI0G30/HNOMY11Qi4qq0pc61Epayf5sHx4Eg2djyb/kY0LUEZrt/jXQNWGfnxSsN
t2mtqkX0Pf+socYWbqk8KujKjP2WJebn9vYzyCeGP/RxZC6JwDf+cWvTL4tbWeza
0e8IqhK4a06W+qKz8zJoiMLcNxNAvUsHLMV5whTp7cMCJ1g9/ekAxcVQDqIvu39y
ZKcnPFo6wfr1Drc1bPqdVJAHfPuqSm6RBKUjBCvFl3+mamb/zE+ZfNViCOgO2XnH
VD6K2poOIpKJ7t1vhONuE9RIyWY2qAsJlG2hemT8TFIOq0w5mu0qwri/oXb4WUFP
VGbTfx7vh9LeBosyEOZ2oTide2gkqX+fr7Slrznqb97NADDtHlwx0Woj/FP5Mz0i
wrOr7FdFyyRkrHvmM4mvW5jQKOcamHX/P3875Wx8CX86ylFMWxVDm8bTwQzy/BmY
8N7M51V6+9vNo8UQr7bA0HRIpyXoFx57RqULJ8BG2aLLJkNMpclXv+a0iR2fVvlj
lk4qpsDuybdheUH9nATcv9jvhv4I3+ui3f1IGM4ksVZyztC8zSAm7mW4QXTGd6wi
rd6fWmqD2bqgmWAvjjUIoU2weF55zofA/2xAmRqzD00cGBolwVwzxEzszMY8TOHV
5dC603rB/dVeMrZw0/awGExPK/ETyQU6rMqrCwMlAquDfPCHNUQT/ogZF9203+Vz
/k8Klk9aJb/tGlCA135ScE/Xicj1gNSsfBvutTuGltjhQlR99AqX5kBjVhSWVxAq
89mYmgEYcOIcpbd6W0q+VqBFhMrl6MQ9VYsivPhNJebd7ZCRbe7WTFk2yBT2bLWq
d1KB7SrdPmJW5Tjyz9BOQWOPI+L4NXakFe1yjg/B/xvgo8xHdz92Tx7cs843AVWw
1mRvYibpJdGPFNhtw4pYTiZ9yqjK6XoGvo59ecLhcxQlTS0bDRPw4TStooFQK6v4
MxtffXxzsS+3fdUJuBYYBI0gl8Bw9dawbNPf4kZTOzdWHMXv9xIvQPaAPi2sRWTd
dF4LSwVJHvRe7Vhf9RCwpAwss3IcfnXCe4PBhmPxGHNvMdm5/1AgZBuuRfYm0m34
hO910zWuzKKVImikDpq0BogqTjdOpaBMGYEIMgqsee53gF5Aa5V0BNmAHBRZBaIM
mSpwWH/yJZ7as7+ot85nhHR/SF/4DRfaKtJTJ539qbYOmk8TmFKUit8tGAdINqhX
QKiQXmJI8CNDdgj+C0DXQWOaZ//wv2sc5W9b70wdDHEkJMGEOlIUetR4ntODCPUQ
eis/hFj+pDzywn3Uw1ilW9V09F4O/priZ4eOHDbrC8V6wXTlyPeLm5IK4oewYvpo
KgMTjxfo5bKibSOfp+tDOMQBEJ5tqo1XStFGKPOkGLuCVDFF4916sE9bOzlHyrHK
w2OVUGiAZbme+ZOFh7isDH4wb+49tTFaw6bukWRP1o425HNsFtEypWPuo86WRwT+
2cJ77lHNq4GPUeeU5QiWvkh2zmFlK04AQoLXQn/skGQYyOk4+Vq3bIIxmHhMHPtQ
o7HWosyitkKlQkOearf88D3v/FGGjHmgtHkBPDPBzUsn/ka1u0CogAoxToODbvQu
/lEFm1Q8bWNNT0+O0/JHKmU5e3fgkO89MGemCquNjZiWHKEdTYJK8OwuLBJgap8p
vFatTh+mVW1tgrf2QwzC7WS1nm5GwZUcwLh6L7eyyX0cnOfaAesNpYmcVh6NME2g
gSDbQrVLEaZ6DqMwA6AiXYitA0gjub/CYT29wUM80tEzHMdV6XhjL6uftEZqhGKa
q36qX2dIaEajKz1bNFpDeYbeuvoR5WzR6A2i0lbhiY353u7JUXJQoj+oYZEaR4UP
G5OLMfdkrYOdNv22uqiwI7jG63nEMuXyURqpGmxyPlYsdXLOCCrD+7WUMfZqZjqU
VYvKf8zMQxpWi5GofHYwju8WHT12ZxktvFbAHhR67GYQ0YECIfMSeu+UKlckmp+5
xqweSntFlDLqFVrAJohCTlPXiwMmnrygsHotp8KfgSY=
//pragma protect end_data_block
//pragma protect digest_block
ipETLYa/dJtzB/57nRX0rpYwLK8=
//pragma protect end_digest_block
//pragma protect end_protected
