// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
jo7VSBcWNqrwyz/J6q8oEcSBcldlXrdeVG9G7FB4SmJHvTwAbnUq7w3nqt1QsxH3uoP6j7hCSssh
oLuDaHgXCkdNkuyTrzR/kONs+BvZXomU6lmevb7tM2SovUxVtm0auFuJkI7XF1+Ui/NHBTsjwsav
KaorodEY+iFSw3yL0M0G1TEDt4YyBo+tc4ULOvrfL3dgGkOIJn+FFeLsjbAyOE+pyYmJq3vm7/jJ
q5vGlCBMR7Ht+79AsbpyCtswlyPoCUd03hOV6NNKR5W3uoSaRfjb1trVfjTpycKMbZ48jv10cTle
b/1qSyQZTsvFC/eVLlvaYJARlQ+6zP/69QV3KQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
8/7AGcTUaNDSehQtrM5haxttz9XUyVIbG54HH27hO1+S2mOYQjrRXVVdg/+BUAcGea5aNCUi7FFS
l5YW76MQMf1oKYRFWjjdqxViALb9CZELGmMlQdAisqJPix0Rb/b/Ds23j9v2qVSfCFSE5lYdHq6s
4KJmfy5o13v6GDB7aJUpPM1YtTsgtUjFhtS5UF3whrci6guWniZcwxpq8O+JjWZphGRnzfROODW2
rw4asyDn9XOnds5mWXTirOGIVRrp/NpqX1UK7P5LHfpnBEuI4PQiETBVubFzRPMsz+c9I5Whvjfm
y/cN5/hdXAEKDb1UcrqHE9d8jx5YchOtuOUnSjJOxx5FS9U6t5AtXjFRyN0EMIPWOvhdqPPgxviC
7UCvjWZbhmmx2qsCtA7O+sEybvlGnFldmd+BFy9tEET/HX1Bkspr9quVELy87VlOJaY7v7p/lL3G
OI0r2JS7DKYk8iNI3w00himThD0ljEwJNlXZPcGsPUUphKFcGMbjrfB95IjLlmruHjud/Xv1oUj9
0s61XW6304U9NiVDwbxIqUJcr45KYk6ojlI25nL53t0N+IDl3bu3sS1Kp2Uvpz991w4GZ2e15Jck
qNv5fdVtb8jw/uWmLjU+c+HI4PI0mvM3HDQNNCFSxVBTBqHNJGX2BUxh3Kk5pJ3QOiCBq6+L3s1d
VreB1WAma0yNHZ/Ey736b7IePxJ/iukGKoVMNV/w/4usEVvQ5Ja6FIXnDs4u/0iv66FBJgE9wymb
QUb0mTwdRgKuEusQcUKTrmaTDxDayBNtcMCD4Hi1mQ8meN8qdsPyc+NTTj6xA6mC6OXaUxmvazfM
ttTfm/C9hhghankEQ4wIJcSTJ+FeX8g804b5BzWo+y2cdg7MgUXejsE01LL2xrCiB9CtCy5lzGtJ
s0nCFCgJLg7m6an4QWH351SQNMA4n8PTsiP0OoAj50rhOcFO13ei+wAHoWf0jXNPYWeQ147aF2JM
k/8KbIFVf86fONWUvPkQ14DkdgvciUAnmtXRfBc9nVfT7HHFcdno81tm8d8ugw215VWCd0LfuFGT
NantPU+034pwfClobAeIRSOFhdciIsMSG1EI2ExKD4GVlpGQSOcw4jmqsnWFJQmnco6d8aEZ3/8b
pqCb7Xo8abZ/YvFMzZB2+yZV0P0HtmvqzIrl70nV0waYi61TCwf9tgT9+SuwE80WkC879Go1gp/1
nj3eWMuS8jYftY9+9j0JqNtiAqKua5G4dm9a/79/Hr+pP5ghpNxytRQdUjo/+7vVRZudTF74Yrj9
BLbSVnAq0rWrdns6ab27fs/MOnwj6UgbdL8qP3JVKNwx0cUT4fE1rXXw0FFkEHca+URanBgNKyLu
bT7PLGgL/zTy0dWyPxeQJKTv6mNE9+VJPag3NGCom4TpRZKNowxSIP3Ggzwl2Pa1OL7PKkE8Qypr
zXuwXm/dmGFzjJGnl1RmwrbwR1mGFbuM46AMchcr2tfJQ9PWMEW9XurelEMvfNomnPwHI2VK6tPf
0M/rdXPLMyvgeh1vCQi4uBo3xe13l9ZAq0MErUjjgR3ka/wyaHQjMxjPwTXtHHJaosU/Boe2YfcW
qi3VknavGCqFaWtMFYZIhSzX9r+2tZFKS86t/2+ncYyzLe6fV2vKD1oboJTocqjo6mVxX76U8pA1
ntVUdZR9Ti57A0eVc1k5rD0H8NcBzZfNeKiM04bZtOaAoW7+eD39jDJyrFk8OtUbld/XHU7HrZzE
QfkWkA55TVQy8EYCheUpJOE9ZvaTutmFbcoqFmMGHGbzbFwDbZ7PqULiz33fm7nQsBQ/KYH9sUGx
nXc000Pf33mj8Fpsc9SsqBC/cZIkACY4Geh8rVqaKIgrTOWp85u8P58dHE1N+Gn5lLBtnOM0xwpr
n8l02JfgzXtDl+atpt2XCHUHT9Ok2gS4mgRGGqJxCiIEJVw1JI0lTpdVkd7/6MLxUj9LCei9+ZPl
z1n8ciLAVQwCNSkLTs/U54ocz4PsCUSrSnWk3cwncFquIN1Ou1RqsSz6t7P+uXniOmlybtL3QYte
gBNhSdcPKnRaHQjxFuSYxQdrNBGaK+ykOzn0kCi/XQD9mXpyIzffNKcG3Ee6Xc1tiyIyVdEJYLxZ
/TonrLrLw8JGhlpxEwMZGHilLRlMXfN1T+RULXJqJo/bs4Zn7GUdJvX+30bBYfc7UtJNnNrrpoD5
ocm9PJtHeYu+VrUuNIt2+rc5LBvKDhuPB/PSlYuYTqVfohnpanE0tZ7vdI/pB28S/wpfGtjhsIZk
2Yru8oXfvrEibh5j49motK/9xxTX9/Sh+ObqxOXh58w2ohEpRaPPAMxc3Sq0Cf/d5mN+Llckrk6q
jIKtAwuYgc6Tbq/e7tDO1OJXbfjAW+eE8ACw/JfGOVFof+WKy22RSOVYWgBO5OlyxJKYGi+tAUIy
HKVL5d2MBno7FxPwit4mYHdcCwN4T3dOBDg0xglQRsJlVNinTwJvSGex5lIMhs7/W/lzWG7bJsn8
ThQNRpSovZF691L2M3lmGqfcEhyvckK3VfTC6l6y20A0tR/Jdw7jLbJj3GCIZzLzo3DhDO2cgq06
G0PwGbP+dSUbAfnkDzWhpIDWWjcbyvsTAye11dIlx+Uz6nH5cuaHJ1Pb0Fv6MPxguq8F2i7IToa6
v4AmlV86C4yBkyVFNrYKNQkiMMXWnLzAPJaU8GFf3Yw7uGwXcY0P9ROg4RhnuD1vq5yugcY1+Nhf
ikEz8RirsAlEy8PFL4utt3P4tIwHdJjToDq67jVomP5mHy3XoT58nJwXa4sqTU2vMjE5LZ6i19Gy
vu0BJtEbDK0CryincGbzEdZplEIw5QI4kfanyjL1MYokOtAA+Gs+yho2Yo0o/cMYsJMmnZXI4K4t
ekFLihw6/wlgy7BID7sov6qDyvCNEfCxpimhI68aJaHY5AwXGNUM0cmfKy+8YbAxGbcrAHhNWoAu
XhXTmoTohqx9lHT0NT+Jx82zOqJyBAZluMnSiz7k7WmfEurrXVZ/YltjaPUnq/8VHTUwU47Dha3Q
5KKU4n0m8HtU8p/2r/FLukeKEGOMzo6/H5Ph9/dYm81NMVQ/IL87ARPxGNPHz/TCgZx6MHyCX7R2
onathVcx5sprkYAr7fHeM2jCmyQ62WEqGnvbpzwQUITOdEkTBbAhxXW9f8T0u/Szlgb8f13UJtEM
6Zg0AG2TSBskIpsaWZ4iFuffp2b2jbf1TOfr2efeUKyC56a36I0bdimovH/9h6zupLB65AYjFs8n
PD5+TxsvErriAEN2Hzjy1wYsLpm0iWSLeJ4ev/YiUABfmmIh+Hzosw+clh05udNkn5Bqxra6jKWx
lR51gdmH3RO1fEZPC18lITWWEucuNJ45sbGcB+ycWWERVbsJihJnyMrmPsVWe0GEP15WIh/rKb8O
Tcr0aXRQxnD2XpBGXX4PlnqfM9jzSZ9QOzqzOFhaO/kLp13G+8yygZb8F36xj59EwqMuk1LdtJss
gc4MH17wHP9T3GgEqaLp5+y5an9ffTjjfArFvW7MoG3hF+SWUO6VJ4V80aM/iUZJxwqh9XTMadIk
TgU8PLkdp70yST7kivgS719Hyqp2Y5paC7KzdpSbxfdgnjTMaSbEX7qlI0BNA3qbWvFBkOIQPudD
KBa7NTJW5nf1JHlzztlZ+OkeWPSFaJldHPA+Y3AMLrpzeta4tkBntaENNCrgdNYwZ/06DF4Npi00
sWjDubzGnJUdU9d2PgQcNY3f/o4KKLGFk2dnHq7S8IsHEWAMwLMUXa3fJE7Kqf6EA/eHcA0ocKec
K+uxQNqTORahuwoHW7am35Fx8YVoUCxIPwj02RiulYUIwMz5c4gSjdG2kV4+f3a48ga4wrOXj8y4
vY5mdkLQHh+xvZCPnXikahISQBmEW81qzXox+MVbLA2iGc3Gs6j63KkJSARp8IorKbbIcj4SMQZA
0E4AVG9T0bqB+82WFcnstur1u/FXikBDmCkems9M/SFyW0qTz5ulof2bwIuCN6EUDmRjYeTPWD8g
jkjrOlBSaSSzdNQyubGFo0aCKYPpVtIm+fyK53S7PXpSLY+01n7rwLipIQw6APdYZRPS0wUlooiK
D8FU++fCrZEbPxJGFrvCxbjJHY4AEWPYrFmr8pq1a8u3v1c4AMnuesdaN4j7kWroyxZDhuztgiJz
AXl1uOJ2X/6iv3YgnZAKTWrHgQvg0JBtDhBGup6npbrSmjEhlyTxrHYmYRZ+RM/nvjdah/MSrODa
JIFyZ7HKPQt7VhL+9owIfh/za6m7I//ooM+xIwucSZK/obLA7k4mkfCPca+Z26m3iCQJkw3Y0JcC
hXPZGeYyIGSXAEMa15o+tZumz0GoMangsCbAg3+HC/xly6f2cweDLUYkZwTKQp7FyTPaXdMpAVIG
4/ZlpWEfntyXoi41SarGtoyuLItxhztWIFT4iEmqSW2K17a/Y2SuChq9yjW/+66qufBdhcwqFNUM
9qhZ6pTr4KOIjy+zqSSVDO/0w2udsk+JSErzew7qzVNkWvOVUsWLmHcP7IPK8aWR71fHPKpQw2KY
/UBrWBiPy8pQK5kruuSt7Ve4hc/5sBaQHuq8L1l6ukcvKZrNj3H3tC50mqlmy+iKxC5QYCc58MX/
l+V/9oD0OTIlzvWmVxo7RWaeUBNzrQu24CdZ+CFRRtF7N6BVPZokleBrpcQN9acp0U6mnfkE9JlN
0vV70VpB4DU6rpipeo3cclLTXsGgb9uSjRsSPMCGyi1Z5aaKHuACPGMSitjETnM/oR/PhzrgXG1C
yWHOLIRR3aW9sgr69enc2R2iVFM6Y4Ld2rYlCX8hfjp9PvJe42jTCaQjVOQPtGfrdc1SP+wEVMRm
MYwjtw2/FCPt/LL//uX5XRmpBzZlWHCouPhqzDUHZQ/gPT3ng3SrEllY8SeeeXhtd3qVGVIF2tMY
vXEfPNNF+LLvnEn4ZBpv510j2bVM4QJOb+UcRDt7INpkCHEb9ANGrGFt7tfgl684bwsspzmzpbxM
kDxrBS2+t8oleXCcPnNNQibmbLinorYB7+TChdT6mcxRM/3Tpjon3ko08JrZ1seOTkfXcUunzvQ+
7FarOhptVJW9QhxeuWLeMjg+IwSGb9oV2I+1C3ZZppSLZac97toH0s+EKnm5XZli4MD1ovt5ktFX
4AeK6SnLXCmplvJt/SbISjPL9M4it3lad5V47JoORJw8issCNKs2Yt4hf+D+ZDjpP4pv/wMHlyhu
1niAqIG/kn6HydgpSVyWUO3HZYMoZ1gHuuouHUVs6rrGNXmQn23lTC2Z2QFjaMdFYyRLjz/yW4Ar
cSI+HGOpLmcdD93hYUvhohsPnlNskK5uW49QMxpVwe/d9vBoldVxkET0NCGcoIoDvc/980yU0zid
3JgAZ9IR2Z6rJFGyU4Txdc3V1rHpg9fzzXU7FN8p4ijba45m9z4OSuVIEBn7SbqdiADQqmQlVi3N
JN7N3UbmYkdXBs2CAqbdZbgK0KtPEmzeTOJ+rM/pbbQDX6bCZgFZo3F42dVxIAxYTFHhdBvXRlDc
hf9OxmU6lbBxkePpm5cSdOAV5P7JYXnBDi0uLsFxy+wllMg2YT8NF2+8R0oe3AVe1Ezi8SxywVCz
OwLwJB6vlKzeYSbcvypIDWR5m53CmBt1dJE0Z9HwfT6JQ4LPGXoCuKax9+8+dnTOQiGjsbI6cKFt
NCW9IQPHEP59JQkiJkv/miqWOv0Js02MpRX9RETEn8Wt7M2pq4JPonsLDOxZSmj90lA6qpQ4vHAw
JK3vmclpfz5RnAb6q9qhWxu74Cx0E2SQstx6Kwhm42x+K+0Hu0W6m7xpU6/f7Bh9e5EX9D1OpPP2
Mc7As4Zc7eDwHU4sVSZqpJSq40sRuV1u2xpoSChCGgcQN0djap4CpmE8J6saag9C5jdyiB3MXNXl
snJQoMwEoDDqGjCgitEsGbwi5xDctKaLc3tFfPareQp/unYiNJJYME2DcAZykpzv3MTu2pYm/eHB
8jubDduk9dxCYto7/P+bSMwj8JWC6ozF9pZmbkB6mpkwj8G+HHivqGCGV/DyTsF6VLcJZPO3AI1R
EOO2CVlgPv6JV5qVmASlvVdA67A5fC5cOsvqk2xubZGd0MfZiEKcBqVCK2mWOYPoTKG0RtN6Jjg/
XbK7uYmlJW4JP5DKt/RM3UCjsNBo1avIQUHd3jP22aWAKxEmIpmHAmIc3/spGRQqb8T1sufi/xqq
H4aSS4nAZT8LRr1t8LIx52yyUWucjqAdk1NlnoZGU5genionvIYrSy9mzIP6r/x+4i30ALFoEG6t
4PgQUa+ot+KP4vkPzx9GJ4vGvvzW1zIWFGlNHRqPzFMbkUuua0oBSEwDFGdg3wSMiBD7NZLtgX7N
p4CFt9dPmvoru0Eru22mzqG0QVEoOrHZqaD0KyIaXsZQFBydbJtS9oanZFXgdTbwboUrX+Xi/4/U
/fv7fxmqi0AnAYHGdSyr/Fj/IOuRkApVxW1d8Nkj6RRF1lpZPzMm9MLa4D1HIRJRiHYWorTdhRj1
IRn2u1vtZGrEuXUrhZe5FTwPsAMwxzszcBeSDMMhzJWOjcflkYPeQanz5f6i2qnLZ5RJxO1bq5Co
gfbDVeUKuKitPICaPsM/8w5XDICMGQtgZSR3biyYPujlju4V/9BFHbvF2ZAbws3H2bDObqgx1LW7
N3bchMM+F2hcT7nmAtbnjDslkkw3huu5oozdy0kzCFZDjPGbrxDI94GC3qnwYl/0GtC59A9mkb51
iALW/WsiaWyLzkmeaavZrgJNhnEAkDY95xT1yIRm65Y5G6sOs2z8gamjHXQVXcxJdPDlZNPA4Yim
PShewrXa2cgLnfeKKFJATswAX7SgeUNsC87pJDkN26XebbPKu6MnziWc2Bwme9mcPfc1p7rKhRur
qfulYj1pXAuoQj4FDWRQOGsmngivwzuFelft9FbejbwggvkqkQHqvuFpu3iZiVZkmRU1jYRd4GoD
5NFsUtxioMhMCGitPhUNdzLqlHgCF54ZfFDpMrCKyWMX23asYrep0oWQgGdeK2TfE7MXfEEPw0di
BBvKkvgL/U5WCOyxXGBOWPJaF6QBLxidH7bdNA43PUrQpgZROpeHDCTHvGgNUnscoxEz/8SRnqZt
knYvD891YT14rao0D+1m6++u16WsLX0AUt3eyI1BuPxqHBaF+0DXadBfTGpl24EOYqx7jN+dcJID
/hoO8gVBaZDfp6D0djR/CEk8RaRo1GkFDmc6aHHNMj6fJnimOrhqaCgxCwjm3RFxR2vZoS+Kc/VW
N6WUSiOBrAkWA2vKbAb3D5XBK3nFGi4uBMgt7x/G+0l3lQEjK2Xj8g7gRyyv3BytHcFB2cy0YynH
dZsvTXP40aMXe+AYwehgJ7RY5SFsBD5nAJFdTik33Pt4yg4Olz9xDwMI8swyfgfgy2CtItV9CCXD
U7F0esgV4DhqR0w0ocwtQmcQxTxWaa0e63JSCfblyert6RWjmhUYQdDtfB0TdRkZzzTjoXymZ72v
4Z5xz8NKHROwOWFjA3wnaHSn9NOwLztKeHIFuSybXVYaMy4+sOVQAZxUWK2DgC7f5XRhAq5813Oa
GN/DoHW39y1RIBNbIV0IJS1FKV9jpuVC/5kruTXju2kUEyZe4RFetkKtL1cMFGsAaiK3dW7BE1pT
lzEZ9D1+KtVY/p7az2cyC6kYoF7VtR4sZQP3Qn4n+VGENAS7ZRx/cAiS4CYObJrrouDGvdVWUion
1zi/3xmrRoBfmlZ7qmeoTU47/M4Sho6ShuB+ldn7spn9RX/sPTG6EAFGtUxz20zblNezT08/qy3J
jZLZM3T3fk4Az13JIvWySLZPokqi2viLeLDNZo8cOf4DMuw60OLfVLNsun0yEgDQ10156mLWkC3S
0MS5mTzO3Xim76/i/HOuplKF6BaMA397b4+0k/g/lIQIuaCHo+P1XrGO+XfILYSchaPhcb78K5qa
7tjRbHyMOLxkeXEr8bhv+kmh8zwJHSqakqQX+gXCyhARhTsLGFavMl5AQg+T/Hq59w6vQf8GduHb
M7nthovg5J4Iwde/dZ2k/5Sto0+gFna1ymeNT1CFS1SroxdXNacqZvSkhfZjtSaPXHX8ShvpAq0Q
DMaCubOpBxbBGa2Rl1NcNKijYEc5+q+WMGJyOZ4eIxj/m7pPGjeZOiAO3CsnRRvmf8ycy8bLPSAZ
Bt0HqSga/0J+w92kdu1I5VEDP0KCMuDS9gz0aTGzCsdE92atXadyRqxqGqt0MZGAlrXb4JUj0VKe
4qYQXem8uNCOL8KrItPTbrmf5g0dmUP6TV9QFgagRuashg20mmoX2oOiEqdgemOQZdcPs2h6926Z
c8sORWv+7r1mp+APhpf5uusxETDdYS1NMuk7w8b5bn4pNEP1q4L9d6pFQSEg/oLdwZZvApNYOae9
X93yKyWg67tsPvWX2SHbLx+HIeuZStMi/9hbzGoq+QFw5SEnZTQoydgge3IiQ/EEMWDmt41cctMg
J81IxMv9r+yDk6NL82vHXvaSw4lOLLMMsc3jEQVMyefdZKxiVpZ08Q6E3Us+EywPc2R3UOBnby8T
ZV0i5VEJQKe1RA8JKXvGitVZQO7JTcpR6ZY34ewoPFoDxcQ9HaJxnYDqPDZuiH5G78Gw9oX8ynHV
V5BEb34g1avrKQk5LR2qEENjfV/F2mpvSOozXBJBeerMfGZk9usNClgwkgOABGry+VqUiqcmn38N
U+/ycOLZ1KQMa88OLhpqAU8iCy7Sheyaji9ZHO1FWZ9RbZyztjsTDLLE2F7rXaN5tVI4HRKgOelT
6/4+5/HJ/ANNLu9EEnlnTMETc2ToKmkUsd4/4AQMyCcmHfVxZwvBMvNdSfzpCaPvpWFXBiLoHD6Q
V+UW7TzvQP3TIJzxzNDq8JTIff8xoPagIki3XWbtRkeZJ9NZgYQls15B9pL7I5qAei6qxS2qnigQ
pD6IhAG5wrEcE5zjJ3PqZcgyndOHmKT6Q+rvKL/zKAcwvm1zhycHbIlUGLg0HKvEXjfPF3mMgWuy
XtbFAYii/AXd8HloJMkOWfnCmvpgu/xvfNf2Dc2iV4j4HfBJJWhCHEr+QDrNSM8rP0yesVCu3XJC
SwveKROvehn/83u7Ss4zpqYmgMS+gZ/vkd6U9ZYkYXi+22+TxvW9Np8+WNS9NQ79Cdv2x3FfbAT5
PDyyJaEzo8DBy2IqThmuSbuuKBDdR9CX1n0I/MeorePx/IFqCMMkgU57RoKJQhDl9i/jvLszREYR
jEDjWTFHqTkiLoH28J9bTvoAiZtEp9rTCthE6P3Nc7YHvUWNKnjgjZqjRxxoQwm9Kczwaf0LUdLv
tcSEwzG0CAbkPKzOabhsOz1enDlPIBfiQCsX5UrV9kNbMWPfIgqH2o+s4ZNoOxWQnaKyEJ5NM6tL
JYX+WwFdMUVJQj4euuHmYYdnBJ4PLWJoauSC5XgUJYrAHT00MB/ygiP8v0m51rP0CcOG36AjsRtP
yXL0H+cRh9+nLAiyihuF1cFelSfKDWtB6tDZn6+ZZhJn8WJA2YAg+uulRXwkBbdwmolVf3vPc8Pm
dUVOKYCOedGo+z91CmGHN55tKYlzmfMS31JUYH0NisR+iSc8BU56pw6M+FQsbXRFAoWLXcnQPMsr
aTTggKIx6QMetMXKl6+sr793znzuju/kOwr5O9WJx+4dCx2c+MUWZLohy1ZhdryON3mPmG3DmPCE
axoH/IBL/HS+Ifcb9gi/s32bZyjwhpg7ZMaleBBiavo9xG2o6CaN+vt+0QoeeVpzp6mHDKxWY9pl
I1uTrPnjmwJl8z20ykb0fN79b9L4An2CXiiz3U+/heRVG4RXWG8beKE3t8lP9K/LcqQv2kmlOrqW
G5d4Q+vvoBngR063px/+VBsZOU1QVlRh+CCKrUks81/oHQoWEyhnTlX38ZyFKxAu33nPNitOqtcj
/n90tbxlUcFyc0kIsVspNBlOc3rqfUk8Le9ill6Hy2w9go8mQjzANuK9/sDd2fHxC7zF4ZtAvrsM
iB6dzQQbNaX6l5Uek5Os5Wzf2osfkwZXPSLROQU6EICXztCphQMc4HdCEC6QUwZPfRWOGb7Gugof
0ow7rq4tej47XJZ1Z3KKV1LAhwVdSzG2bW7Sn6x3NaQSZntkpM4rgLrv14F+PF5UdHUB5Z1BWZXD
seM7/GevyyivS+iREQCJ1ZJC1XFcz8GimrmzpyO7JYMc3mUFhzVrztiq0EftdY3iTSDhWWh5x9XF
q58Mi6/YSH7EVrQBHku7aiCjEnMGUS7N7W3IPKBzPLGpbJ1mcHXTRtLdj+VbGsI4WIfFtraUWZ2d
xImdkHG/W5CyozFPTscdTJClS9fyRw98ZpYxRh0TxCCCvvjiv3xlp7r8+m1eJXNaHg7lI/8/Uc+u
s5j+TCRsy7QumBl5G/Ma7mFTJdgnFO4U+IRnr+gPhUYNkAV8/TyII8B2YSKyYPZjQgnl4czn5k16
fJ90UZomSqgE6JdWyStugPswFEY9YJHYBzondwEq2Vdh5N4+HvSuo0ZPSSNfjDizC5nb+p8LwXg9
ij2PUrSU7BgFObdoNxmoEStX+EzGgMo63S1psVndqlYtvfASSK0ZGIwxSYtyJfNBRxy2/h92Cf7y
u1T4HoJSnsa73rOxU/au081bKa1/oAFvOndQQcACOuYqe7BgjNztmyjittlzg+ILiRfk214iPxRe
6bGc65232qSPfq4/qTE8hbfCqaQFDtDW2ppSHN808ufHPeBgNDcMpD73RAJray8TLXxoSktAK8Kg
dkDJkdMO6OsoHJ3RvrfsHUHtIY9JK+0i9oaBtwt55OODnttX/gf1kgd9C0EBkoN4PzBJPbYOduA9
2gMibm03r6DRD4FrXOvQ8zc8MrHRpx9zwu5WcgxDW1NEXI5Vtn94ZI8StYG8XbYP+YI1reUaO8Y/
uOT1mn2tYJ2yDk+kdycVNxU+vYpbUYwA4giDLIV4UFLTpd27948QR6ShrsqbaQRtILcvPcqolWA3
vG+22OxdxkMQFe6vFwfZ3QiXECEVbECDV3AcJtyIenAysmjSohbh1jLpT+TZtqXg8qEFsfJcaART
6D6Kib5Hfo1C7Uz4NFhIls00kOxoVY1sgl7ugGa+A2dZlkXK6AIPzwKpoMCiDoH39rGnq2I6WCHZ
OptQZei5yqRQbgXJLzPOfd2OOHDeQITo7P7jwMc/3sCDPGWEgZ5haTEc2mNxji2ub0jvKqAoDkQJ
EEcU/5xL9JMdpVeAjK59uG3f7XYmAEj6HwRDnNnTP+1WtCw48sMe1nrXfPM92JJs7KoDoDyVs20C
1FjE7pDn9iIWfJVlbkMEK/HwcFdcGfUyXkGg4V9pRwcQbUFtm4MD4FHnnMS/YmViPaCEMF11UjWM
CZbyBXH4LL3c8sf5ljRNiUjQo4Y3LiQZ0SikxIq0xwv5x2hgIBGRi1S1vHuPfTPfYr8MjzHqvZrm
ofWE/DxuAoM17VHdTDq20ujvYHWBF1aaKtO1WuL+pEoulmvVyBsp5KmakKHOOfBpW3UuftXR+cUe
WaZhIct10KvAAKKF/N6VC/hBm7jMus88RnTIo0wju4s3WUt4eDl6AjtZhyGgy7+VB2Hhx30nRwnv
iByhw/v5n6ZzFKm6yeCXeycgnik1wQh02TUZMDK1T52qjqD7NqXaQN02Ofc9VhxB4DjZuKYFSfO9
ZaV511lDt7wrqnRxVb96z7PazSOIv1DV8sKnnPXyhsgqy2G8WPp98Mcjqkue7AfK39nTilAObNF2
IJDpRiumZmJvqQCSl6UjAM00aWFQqNIuaDvCGQAgzBjFznw/TCP5IvoXpPpZvAOX2D5hYbtmxVWh
Ln5QvkiNZU5pcMKo8Pq3SryCX234ND+htG+m3HUYk0La6eusHfxaRSMef8fRMFfUgA8wfTrzLmFN
wSM7o17rUTUgRZntpl3wxrGY0X5W7R+vpd8O8/8msXkHRCOC6sMK01RcazjowBFrnL+Q8wyVBK+O
0RhSD/lcqC+GskI+rOHKXdSMUoqkM4o+k9dhmDMJ3VCdqyhrIDg4jbN3rd6w4VrYOdsanZRm5TnH
jbPZuHjyst1InQxzBYVzTc0K7oS7OxgH8qWXzuMD4U9J/eGv3Hm+2c5Z4qeQJ9As3TVK4cy2yW88
lXhAc6Tn4qRyFUYR2j6fASrJ9pbN0NzTLVGRpIpNaF6P5MLNRpUzof0cMeUT8ruJnBC+nJaq62Rv
5glAfZkIhXWv56PsdDU72QEp0uuC0fS/a5PG+nhFh56Dp6U7j1AWNi7AMFn7FQ+z36QK0rz8wLq5
IIBpXovOoqeunVJUpAJ1pTVCZ/DD20ejn0+BlnVrghtO/oKiXIhchw6v//SMkpOussDQUVaWnkH5
EnaOrGp/IvTuCzXv6ltRQy7prrF3AyLR5J2/PcE2SZudJHjsR6qUIA2uAnrjQP7m0qvs33CESbQ1
SngTpZyWxwpMRJFl5X5tAIfSkA647L1zzWfCAW1WJ7p2D1B/wV5Jr0Wql0pYJbqvXoepgviySgy8
IGTz7NCHgfdnlEpWiEdPexBsS6Xzjx3GAw9BOcttzCGjTVBDjjkr9Eky3Sxt/JqH7BhWf7hyFXOy
1kdvIBjvnQx4MJMpK+qBBpTpfFyKXJf2tONrLcwwKFghs2C7br59G3JskxJWbSxHevKPPn/zBlmV
iAmnHm32m8PDHnGo96N7MWX+G8ILJufgLFlKv0CB4TBebOJMp2ewvn7H/4x1hySiGDANDgHx41nL
7aawV4ZOuLGwsTjhkj8TfCVtMLMttwg3O8/MbJ+Hxhgd/LUVTadWvl4xRHs1xVWX9hN5U/oDHVBx
WKOWg1f6FedByMo/Wj28RlmKbRLTeL+N8eIkT/m9Lf/aP6Xz+NftiLGSpuD1sTMplv0VfoC0rj8F
lrsI+ffpKcEDspBHmWLgaVR0QNrPd9/yB0PbW79DHPRaSW8+SbTDJ97dubZAVaC3YraH5gjmIrCx
KK26c68az+aeAuiqlV4BW0hUgHBxGblxrZNjBkW+6K+2K90uHa8FQNWE80RPZOEauHgJEwhWXgDN
sp2uTxWaSGWfE67JxSfjBHjalFn/vopIW6KkxSSY8DbxQxcJSmf2CervS/uOVL3UcVWu0dmzTHy1
6x0ovMa3WBL9xiWdTU40HG0H0D7oUTgjzJ8SXrEWw2Jiyzmm4wojYy7ZoZwOWSW2pZdum0PyHb0b
BGlY3gRGJy4Nj6MaIDw/nB6AN2Zi5yKkK3QJ33ONtvetxTsY4cA8fHMlh/qAVlcJue38idHI7G57
wfFdUYI8D9DwcoHQh3Gk7yz8lUjuLvaSHXLsiNHllPhN+wBc6wlvGgC53IFnQ20/gFEhIc4XJIVl
Zg7/HWwNM7H8rKVplzZuJRvt/+fj/C9st/vka6utIaNRyhZtNQ21VuD66O8/wgLKWBx35grm4del
uGiU9ih87OVVA2RAj5tTiakUwuzlQ4pOqq1j6y6YC7MeX0gv7oDKPw32PzZmTRwr2hVYbhnFkqGS
p5tGrk6kgm9JlO247y8Ye/gIIhirWJ0BGWVaV2W2a4+BqExdyWReEJjN3ANTMaVhP1iEDsYjG3V1
MU6YKH88mJRZ/gRgrXrFBxy9sRmagA/YwXHf+FpiNIFNosvGE27UqEQyUM5KKDAI+3ZvUk5vWhsL
AjoVEDhaO5+YEohg8P+k6sMfyfhsiV52azIPJHXq/G03S9dVdQlZtX7/9WeprQLwkBGAXeeVEyiB
gW+L1+jijDO0LYQs7ORSuUw40bvLjFWNd/UZHfPSMJMnouH97knVErOIA43WzQ01poplwdCIBugD
3q3FFRL/oOOaX7X1D/fgNOqYerk/66rPGpOOTkxxaO+Sah6vd01nt2n5LEvsx1/683p2Ewl0Hmad
uaoCwYJn8mj2FUiQRuH2y3oIWSU1nGswmKVj3kY1T9YP2IdayiyKE7JKwDr1mTb2J1yVEmTWPIR1
rC4lAtNabIYRctfaC7JOzGkdsc9STKTZGEOoZnCDPFxKlawv0BDEqOe7OFROR3HULmspdkHLvLea
gr2VW0PHbpS7ePIP7XHJNuP2vDUYBtXMsulmDlwweDIpTv3C4T5856pgbiJ2NxL50XmdxGMd9voA
DwQVzC+oJrlTsbRoCJfEg1vxEeIcuSidmomIhYauIX5yQ6WB2I1piuXDLgR0I5n98p7fH6x0MD9K
iNbCkfmbooaHRd/7II3asQFKi5nSED/InqRGageaSqtp/n2EUfyIua+ntvWuAnDDWY8H1ikp7QY6
SionHcRBYcvU0f9WCv+M3EFWmk9DZEBOCW8Ah57w1BfLdnwy+AX/FEl4WOxgYQ9/2Rqje+A2msHK
Tg4MeNbf22eOph43KrRf2mWUFfKg9gjQwGPlnDqAPnO7xF/mSM4Z9fYFyAOV+Gh3yi0b5DbNy9fI
ZShR0pURbvDGcelWkMDC0XYqEO/dOau4iaLJqWGH/xQEUxYkAiLDZpCbNe3c2K5+T9OMBmy3RSrb
cjyevGxR+LHudAOI1fWggIHoI+RZAHPYos8UhYzoAz/EfhUJmv+TZZ5LIwtVtXZocs51iFv2/nEN
sckic8JkM3OrI4YHewqSLTvnnDauWUHdlvlJQzhP79avmgvahVNhPGD0YywN6bWAWpf+IYu9cPMZ
i1rRdTE5plnPgJNznMDYOCVURi55VWEDRtXQ9CDHO8Mps6WrJVbW41tlLP8LXSQFXufFXIlgQrlA
4qk5NnFn3lLtTzbyQ4MFdWN5lulv0FAY4z5TuJ3ayuY5kFeJ7qdaW2DanVwxtwX9NACtGZAlDyvm
hwm+yCadyIPoda582K9Nvbuql4EOs94lnXoRM28MJ9pHbImJS9BPcz/xU9tXwk3WJoFbHNNN5o5V
qVAsVuXufNSj1PC7CBdwWRWYtiiN7Uj74Y7Q1CSFDv2+RuKSCIJYp2+kBfwhORQH7qo63vIxhMmw
Nq126Ies6p4eHgio+c1nMUcjUH8lUKnajnA8om8AxKfrWllre60TPANLUlF1vzU5N+dgR+klW5xd
kWpll8mvJ6cUvmOKUvTFwqDxezWrZBP+qSRcq9k6wBn0/D+nrdBtxnjDRoclqSvvdW/g3qfRpCZ+
3/ec+0nKTrg/80fi1sBdx6mQsywf7Auxkf1Zvm6zU4j80v7eYR1/ZoJ3Vchgy9drzpam+EJmEh9L
yXawXmWeRAoVYyB4L0SJT97INbbXuMpXMvmtcLtuH184ffhaC3WioG+qkz24j3zcxn232vb+gwAz
APWbyfEcCTx7mEcZZJvBzNTwSq10MdgAljn6WoOkG6bKjt7vH9Om2NXY8zhbKYa9kbzmVMxKE30h
sPTm6zDrWva3lMmJFgHFO2vWnd1pkk/LyJCIeylGtwt1EPkP/987W73ory0pzgxqcji+d0AUgZQc
BII+JrvOM8osoTFbU6hF3kcgqWWPArCpJNKM9Z/KNq8mnERt5jWnsr7er6q3jqh60TOKpXOnQlFp
Wzbt7knGyD/NaF3EtpAXv+Pko+JUm6u6cIFyX7or2gmxLV+FPRqAi+uFUIfDjj4lJm6FkF1H+/wR
7SYt+pKLnskldVKIvVkDsmZ4CZl7TKLjoqGJnlo4T8vtnwjRkUmwTWNbFC4QYPX2PMINhf5udgnv
Pj7oEF9xP6zaHoPwN0GFuIHWVTxDw7MXTVxRfffUpQw13yk03Ywc3Ez9eroACKMFL+3yNb1o4SoQ
eUHpJ+7Cp3/njy3dRRdQ+oaouhdblLJoS71FXx6PEFEMk4AxvzYK9FoSA/oaeN1mG4RxQkiTyR83
Y+YaLPKh0lUK7Dp23PX6RkMZJsSpfu8JVIy8LocfHxAVx6l3Lx3evgxubRSM3c3mfYixzzW5H1R8
nDY7XdJbncS1+vCf9PdOHtcnJtfLrppHH/WvmLoVcqSbcDEqw5pUxVF7VPA5Rh9JwsCRBzB8tH8w
W1XCL4D5Dl5HcoGTUfKEHgWzIwifrdYNQ6tuLQiv2N8rbtYFTaErZ7DLvHPhyBIJ0pXh4wuLNxi2
TGD+ZWSIL8Hl/65NRGXy3pcjG+7PhRXCj+yEpTc4o3a016x6FaNYaH44MyjjMoRB3Uad4I5oN7Jc
a6oj04Qy89bVEWkCFn0ae0KuJfLzx5Sc/M/hRUrW8VDuzhALv1XOm7L1vPlD9XLt4r1GTSFSUJs+
BupifFRSpSIyWufaxj6/iAyDdngzIYFJtq0SyKf+j+Z4GdqqTwQ6gfs4MiP1BrIeH4xlKR3VITQr
7Xq8aDc0Wvi1C1YaNAljAAhzxpTh+qDi1kT+6oy/Y8mOZh2OYzG46TkUiBfNntw2HXgXWkROyQP9
XryB6XjXH+GfX1fs9+IX7utb4XfviX+55feJgiPj/2yFrlV3HVSYZLKytBluSllzeQAFf228vWW4
qwofu2c16R2EkJ1OACxPUVkRieYEIMWV7S/QnB9AYHy13Mc6k4OgtdxCZimqxGlENFjAbIlrQJ79
ommWccbetTAWee+vS8nKPfKr+OJ3TtC4OSpnt/PXhSUB2b6+naAEbH99nVlomCYTsF89NP/xay+u
AO+uopVczYWWuZCtucdgqGGDytEak6EzEWnlMXqYdfqc1zNOh+Ep2zzKpKqfi4A1E2bDjDF0UyDD
FxNIWvtWgumUgBpS/FUVwj9jHRB5i3zo0xMnCdCGatEFlcEjG2rN8iyCJiSp15BRSghSSGaRltNf
gfpd48dusQY5yZXz56AbTOlIqHKOdVHeHmWs8UuoekM3QunJXhqr/yIxph5HS8f/eFjq5wJHr1FR
naqngTeZVPXwuz9+NJDxn5EsTNLYUh6E8IW/cDEe5u5h2Unf8QaGPtdT1bsrnRV0P57ryXQRYIRE
fZjHemwEGezulhXjEu5E5GqSX1IWn0zJctrzEp+IcBHJB+2fmMFpn0wDwGjQI1odvpOeCQyrC84l
VsGHdXPQ6ENe/imiptJ3In59GqcGYWf0a1zOJ6FPqYGxyTXpkEeBbIxN8pMT9F3fwHVJGN4Wtcr8
B/bgKG8ibsb3X5VXay3nhbJ7ibOy5k4yfJtbjaH2AG5+jXHiYf+KLCMVbLyDF4FBl0ZF8qX5WpzA
ZW5ojRczpHBE8qGv67T83pKnAWXID5Lew6yP7eXMl1OC/TOtwZxw0cdAwOLkeGqJn87+koWjvMYO
k/bI52csa/02L0xPyjuYhxCQNffGaHwFBH+jczoB9cLei1Iqfx4mC4pBWwjFmHH+58uigkOfH0Ji
FDyXOrwQj5sFMVw/aAbvxFrMUUWvtNSDbqVkI97Kh99EEzk7vZZ3t85jvSlwafjOB25KF/DRwDED
xEffIcBZG+Ou6lA8nZoYn/+qrvvcJ6ZPM8aTQ9idRIMUAxSWk8057fMt93qXvSOrjJD7119YwZ3T
NPNiq86bpHD0K4XooTRHRzJGaCncvdUtf9MM1Cxsh6kULajw7kKYfvbTiSVCCrTvdtHYaPEa+20G
7iIkoAR9ZplzZUrGvwZMllx6kejUJT2hKD5GNlm2PXbusPFBzzimHShLTaBaRzXCHAAAKizgsiFA
pMs3rGmDSEdq5o1Mhp7s2p0mjD81BMtQg2M+veUzyjbG7CMlETUbDnN19QIfvZ4jaysZLQVoQRP5
B0toeFPNs0kTycXju0G+QPCpTkroXsGXAK39tLobvGMJY+IcvOnfgOgs/E8Q/GqDY7jej3DI7gV0
axET8KBU9Mx9f0Mu1cBfT+easyXMi6sbmb5hxgeYGAlJbGUWquSXCYOYwvNfUt/dPMPmSTUWVrdO
aqwK9x1eyzKb+JkZlKtdGScWp/vfyLzWD1N9fkpVzssaMrZpoZSh80aFWXzelWwrktJv96kSz7yJ
3vp3Fj8KOA2dFF56jCYxTpupT57rkIvZudy6yCNsTAjZ+NuzzfhDMGAd3chDi2B+rnwRU+pqYESs
JXVrD/1iQRxJYBL4oC+ANHX+Iq93kn5XZ7gypUqm8Ap9menkqCUZacsp6EfoAeVNzwSQyiX/k92M
dwCIjeXd8ioxD1ADAvupjicNSqQltlM8+nZYzKKHz0uRU9wuyC3b1UqtNokAXTGgceF6Iz/vO4Cb
Nl/6sebNPcp04Ia1fqTwV3Gf0DKhW30jZBJxDKnmmTHkUQBFP6ZuknJ6HjghZ1zuGrAmFV2BDqEo
WwmzXxdV2y0m57UDojbd0goj/irM4yyzRAsYH1yU0Dl4t3n0wlVotEdOAY22w3X/YKF72Fv5kCiI
SeztR7xj6iVYdLIQXx42hj+s/ZOCxONSlaQ5UQ7T14Wrkfe4i+oomt3S+bKZym/40RQnXs/RDy5q
gFIhjpAw8E18FGlzza4y2tBgy4MBNLhD2X6fOzhD1s+vCNsQnO/+6a2nS9CZcuzajyMM6JfX67eK
8HtrUvTPgEmBKfy+sobhdO96ddV22vkJWUQg6b2466LxSiKSBe0O13qGpyppAS2yhIOUHdp36Wtu
4sgHOM2x/ZG93SwQs5mJYJNDim6hstgNzoeEm0wyB+C+OXxbT91pDuurhcMLIzY+/mnxNiEV2+8U
cGg+KtWEhCpqUk3o3FR9v9rzIxzec6benY5QJ3kFfp5ZRU4HCIG0UN4LJ4tVMJtaocQb7s6y72QM
KhmDmi45vX5ZzH8jSoVsHuPifSFyJKMf0/46SjKHJjImgZCcxsTY32XWwG4PfZCTxj/kHgZS6BtO
OG2WDLMKy/fYUWKmlPiIwbFx1r2PPDmVN7zs2hZGYuBDShG3Ktxkqdn/uzH2dHg5RT2sETa86Znq
FutuNPwC0NBxYvP9UPe9hrpmzQOY4sE4TbXcLKPiQ9HLyRmFrQAKSOPm/o2hj2XJKdD/zP7Rcnq+
kZBhmdKcAzFh38AtuUjRcyXl1fM6zX+Y3K2EGrDN49L10sRWDSBjMmLxsA9NbLQ5lSCuf5nQS3Ir
iA0Lc3+9DHOflHkGPVuB4Ba2c12qjN5eYcagItCgNQmpsWHWhx1HmzEZg2Db7H4Vthom7O3y4tHD
2XsxorRSLUmJxvyoo9bOLS7+cO+UG5YRyl1+cBmZ1Pt5B91YBT5x3D/la46WmGF0t1SzmWAByXgr
FvZpu0rKR1dw+X2+G2tVnpKdhV2ZuJVWVY1qBQKX0zqzkR7im2MA9Zbr9P3Rdrnc1z1tXec/k+1T
GnTLekMIKLZGbSEXvkzmKAGl1ZnMWzGPHWxxmo/PyJG4jIoQDNuQvaA9qMM14kXd+U0RtLT+0B7f
GE789D5T+FwoQeD31AGDnlxAPhpfou/iFddV7s2zg9/ei7ARC6CQAj5qRlLEiF1D50QiToNcY2OG
0w2kzI4JTLUZFNFDb1mD5NA+abTQ5QgxrrC2jW2e4BqmshaBCDTko3ZTNX6vN8mkSoYtUxwzFuAX
2mrHwmtGeT6AUgDj0Z2yQWQmrP6uOjtvO/MDlSUGJ8rFXamA0ZTguSvPH6eb3+tdYYyn0oddbnmg
UUwnNDvtdQILRK8MyQtFRCcKpeLQMxe1SBfUTsVWJZPTcPY0CuGYSNo1DLYeBA6GZJgXG6FXXxqo
E+yn7gliG9kMOvmUEHVw5S65B6rarE1JFehoGyX0migzsyOvkU8jCDGhMih13xKKTiBkc1tDB1Mn
Ay2a9N1KY+HW+GPDQOAhPiR5wSezqc1pQeEm/DFAs/P7NRz4S7GNu9vDdHhfYVhDPPBQmKr/Vb+L
XvOl0mZIqSRTNUvAXxdQM0Uhff87nOURKATAapw3LiTdYjZkeFCg9jpCrWaJhgciSo73vtgJdLlG
DxBkbk6PmdWzLNptmBEBCcChC1+ohcL7eYHgmVpf+wKqf1nzkuRL/q7SY5A0k3ojWbVYQoQy49l/
fHwJuXmHAnc/4OE5UN+YwdrAxhCUpmpao6jIeQqesbP71ROkg0MFM2S7DXw2gw/1R1/HmXH7EMTR
BLS2Mh9LMG0uTY6QvHZ0XD6gRvvpuTabry5dymSf2hj4ICroawJCLKktE3qdQH0oHMT1k1DLmvIT
s4qYZiGANLZIluShkG0KtWdzehz6OzUoetTDB+Sws9Qk4j4lLNiJ69Czrl7ohaHObYIzwnXPGfub
wqPnxIcF0OGdp6o7f2o6Rw6zxrblgPTmh9MsJmHO4uV6+F5udVTSoQE7j8ULkwjHthsTTnOa+otI
6bLKuEA5y7tnHqmxq3IZ2c9JCA3VqsT7wBH3wPSjddwZ51z119frgS2QmemYBnySBVAqyGYYhD0J
51cNX9LV0czun25WyT+qeFk7h5Rzj3AdnxKu59ZNcWOsFRJ7jG8NU8kAK68tTq0HrGZhXzlo6kOe
pyVGrlFxmo0aH7WV/28BjUXZmyO7wmIJnZO6XOliUIv9PgSynS3dYz4soTyqSasHlS3TlCLI9at5
VHnYeSInDbknYghiRMzPM3EfVfmgG9aI46hnvpC+BZndeJJc1luUpDAnL9oVCAPhrFU8HNc+unxs
Gz0pPhdPL/0m4OBHw4BJ516sOlLwmP8jypo/e0kz4UzQA3ndCh4F6RMTbqb+0yXGRD3mbc7K+neC
6ajg3lrWTPqDeP+HUSG9OwD4vuMMU+z8s9bJHHDavKoOdo8LMg0Z3kfOiEAiqGLUvHab5O+iFrbd
zFMTd1vodBeZ3wJR9pDwY2UVUIWohb59zu2XNPgZ87aHn0AOBEQ1nHw3Z7XflUqTyUaEID0MplcF
jA26bjA+DxJJATKIUOrQTAOOJBuNzbRJKrIMsMw+DWXeJd1I6Q8Db7vovEGvrCrPtFB3cBw6fHxp
fW6qMqxeY8gOEesKNNRTlrWdbJA5O6+cMdaRf58T1EssYRfJCnB7IKK8/pee5hYM862kuVNEQRI2
0FrE6Nx4Votg8a2dBUGpGeZ+nvDlLnYizaM2rOw3/3sgfOB7KM8KOUQtij/sR6/KEAhtpnHA5PlR
I7gd+SfCy+4Y1yIC5PonKW3gaZaEDH3nfReZESeqESNk0ezj/g+71EiEzdOksGIwBSx+UkhPEhiu
7BmDwywMhSk+It8g7xhVDspbUQT10WiqEs2CGOeQZmCjyqb/7i4dCwMxwc5sTiAGyvnllng3A9mH
Y3NnhxTIxoXlAnN9/4Q1Av5kRfoqJ/e2YRKsQLLVrf6K8R6Fw65jw+U5mZaTnVBs58UGXrJ2sAAX
YaTp/+mfd259rjceEtd9mP9FB1kVeHgM7NORgWzYkds7uEgkfkeo2MSTKDKYlMQV6Fq89jYjwSv8
a04kUzWYrnDYJo9d6tFZxloVKLT31rZD+Hk/PwnY8TxZ9AdyTT2He3UIqQOFY21pngYWfMJFu9lx
SqnwW0T1Yp5Iu9Lwtzf1oEmqvwiXvx58XK0zT/Pn9D0YyuT9Wlp6F7al+W8Ac92ZGszLmjww7U/t
GSeKOqxfeYG+OPs70QuLKvMANJaSTCOjIfoZtcxlsGAyozAtqFk601VNYAa4XGhuKE7BEiDbhseJ
rZb57CFkC6t9Zo51Aihg4beq8p2eyhoCAKUzoaoPttLaYMghWvcRaOF+l7RZOwg2DmylOi0gd+/E
DLOUnelxLQrlISR+3rqetKXb9KRX1bMlwCmXNeQNoKKOIBGtTx8rQ5zhK1sSM2DQNSXN+8j+8Avg
uzUTp+0jfbVvnnHjsY49H4T01alddJ/7REjNCMC0JzcR9QUrQFVWcELLJktRZj9bo6tF7zuOaYGX
sBbe4IK+Cd2y3CeCdbxdqQ2ItAbptmbgEL01eccoqXUfCHd+U1GMmK94NAnrdImxEVmlhR5mrEIK
XGFHoQaGgBZ6hhkg2S0OaZbYEA0ETYyrLO+TRbegLZZyp9fWAChVxAD4YR9gZqYJHxkrLW7AOL/c
NDgVk96ToFbJsW6sAfMsFaL29Jop2et0eiDXRJ4/HzqCBiGdOW/07aQIbfIvRR4/ls9tyw8z4IlD
dHk5xizx/2s2Gg3G0LVtzKmVEBXpEDpyeak5i/LKnOTFMiZcqdOQnlvymrOn4om0XmHja9UUXaur
fsNAjiqROnv6ptBN5jJ8cDG9T6SeCYDxOXRTMyYReOgTsVZkXnHut9aJMM19TxBERqK7jIp7DUu0
5ma6Gbxy1213rN0jbvYaHO3K90BqI01ADRJz1kKGKbff8hhtMvNz+UZeCbJwkZfagE4B43+HQNEF
pvBmg6I8QO4MT/G9NHtFUH/Ec8ENhBC6aV/rpiSowUCpJ54GRPhW3xFw88VSiQY7/IsENAKxp949
+8Cv7uwDgKQCE5Qg/OQYRHSP2HObdinlEKKoiywds9ULQJ+ikiNU3+v2+gCj/K+Wp6+UMFZSjl9z
tpiIn2Ir2ij9SwHZTPWpCIzK4BsJg7O7clPWSFAZBYmsGdBokR1DXhGZ1WhH43nW326eAEv2Hx9E
KtWaUgxNfV1cvHl4n2xPjIkMYWtq7+PPBWUMMUceqWh2raXbZCPffm4h+4D6+p8+IDs+eiWUkd1Z
/4k9L/oS19Wgbh++YHAGRupj5UrtQ/3+7rpZJvwrXG4ZRWt426Z5RC96GjVkagM+wIZQIMj+pMv/
Onrh2P3s47ceSq31RtzAPWfHl1nOApeTRHZTqSuO9lLmsApyL2xhSCe0LX/wtOJDht09vDGcomR2
GQH9fwRIgK5Sp4OfEeI7UWSAmHPN2sU+xB0JvWkT7rVlWLu5PmNzquQDzZvD4jdIf3rMmc5sdsin
RekRqTlRE9h0M75DA1C0PJhN20hzf2/rwHgNaO+yTrjZUCZzG8ZYi0I84wbFR4p89N2FZfI+cRb1
/64QEvpFhKeK9R4N3fm7UB8ayy/EAPNOrfPD2W7aPqS86Jjj80PD/Wt2Z820zQnX/pRqz2MGTKqC
mkPQvEhgKIoSX/6ADIJUdwMiQzcNRdsIfoKO30kpjKDDhLl1W8LP4wfJW1TJJDLtcVia1sR9wWcX
WECgX07f7EQva6/duTPLSCiFTKJuGu/0Fb3pkjnOc788WEO5IChMJ5vSvW3jnNNq9XJbEazl0LvB
6a9OcLlK0ZzWLHRbDDEkpgVAXloPJhzb2quNJW8JFDU7nK3Pt2eVrNwnVqA/9ja/jyo6VEmRLz8t
irhKmFh2ze3jyEb5MVZHXC3z6yjiZn8FW1S0T5anMCtfH5A6pWVhtoWPpbv1wQq00rRJxXvF7VOA
Q4Xhl1LCiOM+ijP7LUKB5RcQkuS+MpsdVPR8r1cJOfJ451XTe8IAN9UVaI1ukonM14OTZR6sz4RU
cUF5QO33mpUGlFyvKkcAm2ggJiPZD7+bAY7wtXjcTsKAAoPfzA6qCDGBJBkvi5e1vK1NIpMkDzQg
LHOa2UZl9RYWklYbVWwjV2ysp7imu9gghxXITrimffF+KixswURDcN6TT2HZwuTq+567/9q6T2zq
0qERPexZFlHfqHhmpivA7TDjXumgoeFcD296UfgDSwkzken36QKuWC4maC2YYM6SFTt/Dn/fcrZ/
fhbtbW2C00m99SbxcV9k5ZAxrI8qqswYvpL0lSn1PreiYNP4gEsQE8R4/aWvGTbIErW2gtpZqYwv
gxB0Vhuoj1SIFeyahA/5Cb5rbSJ7V/qEuvjoeiAPWgsPGmgjmvjp1ZlfPmi+gUvcl7chDpk5RGuu
RhUayK2CkovYAqzfc9CrwUUa9fYeWJEXDKrZTucCHnTpstCxqbHS5WGo+S1FQXZ42TaYtDuc+78C
SSB39cTkJAr/GvbvvyCGbpam4+dMa2YeKuB16f7ZbqpJP2PpFmnCiWUFJDdZw6HR1v6Dj1gG7eCY
AuuhUfl9QyQDE7SKiAOUnf+pP9U38bzJbykw7OfAQm1jrD6LUJvo19CjCsypqDxl5u75ptCCoSDB
E1TDpFFvcCuv/8QVqU1/YRo7XV4aPZdLXlkoC1XQS0Wo9PJHXyUFl7MzXkEQiWg4BwO5aHuOUtwJ
InE3LjBASrUbkmmzxebWEBA0pO33AMyDS2ewuA3j3kb2mUNQC+gVVJmzpXTMxyzElFCSN+Up4ybC
s+qSwlCMFoGQHUTwOukz915X9/33vcbtD1BoaNrXS0xYL6LnIIAOkWZYJkdfWs8ylJ6CximBwntW
ltLcpYRFVsP7alZS0l3OTszI2EgeMpPoERU1GelTWAAoYxqBjJCOUuEJnZMGLBjWgfk07UeM1bgk
YmpsRm7ckpFkJ7oWA7bmld/yC4LOPW0dfoaJSOfKB5SK8NdUftO+qQwS/JP1UPPB1JQ106QL5ltm
Hl72UNdpu+1vrRK5DxAd1CPXt7x3gOUZ8BXC4y34w5mzKTM+ojRuYt94EhvVCjgCCgNdbsX/4vHc
pxdVouX1IC4dNq0tdk1Io/MYpSYJ8WEgHuzzMb5o2LdAQq0sZVFKLPJiM8EEfvCEhpgNKnvinPud
oMhvcPOGd+YLHlq3C6EZAMfV7GRjWO6f41SJ+LQRGqs0IO5FazcG6fU22Iw1FHXN8ChQ+k4ySBVd
xVtB+QiBxvj555bQqkym5+L+oTRRsETmJEyKrcwGby+uFsZHnOoEu5Cgj1EJLaWyF3tr7EgO5eEa
tptqNKvo27uMW2b3JIWpFWCWI8q8MOy20NZcpeL6++Fw4BS1YDNWiEV2nx019JwRVeV7bccWrE+h
/UMNIme5DfuTwwHv9pEQRHuMvdo+IwxRhqteRbDsxE54bw7j2TZqpjyPb0z6KmygsMP04g2c+LlP
FVdB4mUakKnN9IA6KpIcuBL/m3GOHxRpl86Ec/5rfNnj2gp8wKIuSkwEY4nClYM9HAtAcYDhYpmY
1viQ55OGoYMqHzQlqvg3yVgNXhPAEHwu1SttGW8FKjVO7GJ52zBFEklQOISuyIHQWrhgGYrOwAG+
qtQXoHGZUXoou2mBqVb77zZUGrTo6lbOBhxRHamTbLhQ01KLS9W8aPNfU9DV2HOaga9+iDFIMsX2
kFhYngZ+q0GAGSbPxsJeIBzTFuV0ThO4fah6ITa+hE+QmklEsqmUSPvePZLYfd8Ig/raOWNCF8PW
zNrXlVZrq3Ij+cTSryHp0afFCk+XfGoiCfImIjX/Lnl3O/bpvV42e/Fzwb3RCxwlqoRads0xa5eQ
Y7hLpXt5euGbRp8ylW5Agwfovvt9cj/XAYaSLIhDtvr5yOaOzge3EdcableNJB1EhqZoQq69uPi8
m5v9m2JVVBDJZ7jhai3D5cz3Cf4GulLo00n4ggdTVm96bWaYhq/Y0sI/4mSOZ3l3LBcS0B5pNQLh
NU9Tl0A31rq4zw3Pi8K3B55QsF7X4sHGvCkJPn80jPrdc5SBILHULI6UkAD9c2pfXkDeBsmvfIYQ
MJ5z18IAgbtR5yF29X3broj9HUEWNnKBlIiSNKXXIyZQfUaGagJWyIqothnJQSg9B4Dk5EcUIUtb
a1/jlQQU8odIfpv+4fmNp3nXKFOc9vi9fwIMcx1G0SHWEv3Hz1RLMV8Aw4W6o4JKTOrAV7iaXzpk
f/7F8bAlp9Okorbu1D/E9k3+gdSO02QfKfkjdCvdReQ/RivrlMjfNOyu2vDt/ZULjTwhTH8xg8MN
KRg1ii863PreOW2yz7QADcYA5duaTVLAuaT9ugvGErBFmGY2VnHVSK5JVxwKRnscYgRd4cnFbHFL
roWUYYnrEyOmRwytcvC6iFJ80SR8johq5HML04AlM4FB14V6GZGaK011jQdD2obRWWv52i6B74PE
XWRzcciHp9EpfEtFfLS74DlgiYfwxOWnRKZz4ddhJ2OhQt3VKbAWiImQAhKWNvxZweES+Ybr9gfX
3tbBks1hQeJCiuMOihIiIpiUx7sgDNfP6xZd+4HaI18EN1sURPjTPMhi67Tz9pv4AIVCzDDnFPRJ
fCtoniKn2RO/w2JJ6S2Ypr4XUjLP0c/0o+HrsGpwQEBc28Gd5Ord+A7AS3AVcnPlCi7k4EQEf/l7
zwpwRaUfNyoeKnS93ezLVEW4JtL4/6zuY5McO8+gk59jdniOe3nqRDXR0USm78uICrUm1bGvWImJ
Wj0LacmNF6OMQFKP5GhmaurokA0M92+BxAzANvC7xbiTlqHIQ3uif5cwiSb1f4ffbifLKMl0JYa0
Rtp2IhI8UlFEQTWJNnL8TtCyqQ1aoDF67aa8EATuhJNI4InwjKWMq8QI83fUuWVIqGpipCPjY8zh
qH4cLVxhR/botD56jWv4o1yodIcTpt6hVwhs530BqtSb9lYPthaOKb9AbwCeDd62fIbJvKE7kQgo
mGF/lHOkUBNFMYyUQaM7V7DkuyT8bPZ/er1E9RiC6h1Pp4118hMhWal9H2NDIzGmqw1Ya8qaUC/0
ypI3VnrUCVnewkyZVDuUcNaGEmbT+FOQn4QxRWtLmkBnFmEgaTGrpI3ZUE1uQdCuZtupTUHmaod3
QT+ithUYD64Ww//r6D9Xc47Kd/0vT8soVT0YA8BADCj3j/lzEBCoJvdrIwBB4dediGiZ+7biMAzi
Bamxg91zTWROehlYnS7VFap+Diz7Gy7aJMn/XwerK9bUMfhYu85UGo6GyJgjnE5xV3Loray3fmxc
upbi2gpih9zrwB66cWfQT0NTEDFoCWuZV7A9IwKMYztv1kgaQ4yxi3l38CrrvkVwP2YtdaI9yVLT
e5bBVDZ5mqD+qWphrViPuECk53ZJ5yFl0qsYFW3rQ07ZPaPcqbUcKI8xIFsnbLZEkb7wINCDzyz7
8FbQCIEpjr4gbs8q/dYNo7JH7xCk61M/G9Kn/J28MXRc53em1SkKHMpLnKK/EMR44MdYy3n9ipJ1
IGMJyAhmNAAqjJo3AIMMwx8tdZIYJH6IPKEBN2+Zr1SGv/iwywNAOwshuSCF2ONPRj9HJhDj/cMG
vZfdVV7w0B6L1fC/Da3uFFRjeG4DbUKzS56oztkcsa7NL0OD4Esr2cdi2RvbR2z4Ly3CdUzqckBn
vZXuVPew5NZx2qU+PIwVZq7OGDrYhxBG8//nZctBdXRiBvcS/IPv5H7Cb877rUfdMQgHlvjfrjAt
8rnWPXvDa23FBDD5Gpt4lMWFapStPGXrFKr95k3BfRrwg7eFn4jBYssNp8uNAAm74vuomZmA5lh3
xwQHQxkshwrN4Qnhpi3QBhGEtGM1tlRb4u4dpGZm22XVukRwwXV69Oucn3faO1LizKCPuFM/xS35
aF9KSGj/T5igLTik6VxA4VRfTwaSoFc4mRJdaJiwa9EdxPj78S9iW3vtaAsWFmlnc41RGtbw+oqO
LLBiBvLKY+7PfnUi2oEQL9Rh+9jOWJ5FNJab+NgW4P2yCEfjkUVVEMZNDrzO54HltXXKoxlogQfI
akYql+Gi21WhKsBPFPfaHhR5IP/pPv/RfX+kxOb+lHxS1ZbnyezK8EAFkrIbLv8SJq5Wv1lHsp3n
P7yQGYdEMXjZm9os4us8HESiiT/LS+/zr4HWfMjd44RxKcUvDfvpIN7ZzWzxMyZXROo49shfQ1bz
+3cHkQKKuOfvLgLnTKRPHCmRvpA7rYXXv0+NEQN5LKUiOVxh75hNEJmpGkv95jq5G68ClphtzEut
FkUs5BXwNjEl/ygjJo/h87m/dCJLczp8tqkpG0eg7Q3jULqYaGJDdhbCB/KfFMxnV4nOJTCwNsm4
Ry+2Ykz7AhtYzwZ2JBNLeGCP6AqOoxVpskSbZ+RGpm638fNwCGTSlB9kQZa1o+OSIRX8LqwjErP7
lSmBKtcsFX/1ftpAkwRc2CCLNoQ9TZGsOL2HNo7yHAfBSTUAawo3CnzvOBppkn6YMDcJhz6uPGTd
L2qQAFuyyvYfIz+ATQwDfeK7HwNfpM4iJli9yE00L+6baWhg
`pragma protect end_protected
