// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
FO4FwZ04RkZrGJn2bk4kv8jPcmC3aOP28M99RKYO7aCuG08RsLte8V3HNlawRToQYr0Jtk/gDn1y
178sXv9GTy4RjeKiVBKG8HQyeMbZnaXpF8RDDReZn8ZYi5h9DLCo70P7kGkzPbW7A76qzpXZ+2VA
m4bhhXRqU071LuBvEic7r4T8dQPEGJMXkfZuAM9VkaG06mLAUJdN1PMv7EgLqIUBY0KS9WKduR4a
MxvU0/5uB97hWo5ykf6OBQZkSD8+8ZEjj9z93TDbADa+vhLfmSgGVb+h7F9S6dlmncdgUEUelkvM
OWh5ofwjhj+smhEri+VM+ckAdEd42WTTPcpGow==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
sIu5uRqiLQJ2tjWG0g05C9QnSiJecWY0RRhlro7pA3+gCLD2fXHDUov2IdxZenO9QAeiSiIiTMp5
cFbTkZf+LO4QMqFdbZVqCF+cS9vGacuy5crO7H+r8NOQBZ1gFMIHAgM0rdas5279GaHy8DG42G2+
nbYQggDSA6VGmE7M1jKU0XRwgYrXgzVzfHG1p3V7BaBDAdBlBpGPVjOT0dkfl3YigJc4IECJxyTZ
U7xi8dI2zufXKyrrazU3HOZEIHuvdyPhrO0Mho9vPTbZCPJvl1vjNGF38cpeVCoxaeA1gUuEeo8Z
XsW4ovGhj+0S4OAYhhNW+GbiE5h7YsobS+V0cWaoQjEySIU+zw+Ei/L5pR9mWPi7ECOB+PwguYFU
eV5aYSGX7ZOXObdSvgKNQv0nhSdUdfgJZ6QaxTH0Oy9HeBDK6VxMedGZ8C35qmw6Zh5qzoj1piOf
/gfYoTvy6JG6Ue3//q5x+PH2XEhVAXZuYkLoBiPtjyAX/MI/RCzOV0KFZqgwADeRY0eeyVHLgeeF
ET6DBK3jeQ12EuHfOPe1wFlyqDfRdjQd8vNCwe+hr3k1VXKKKUMJ5KMH6GM6FDQ2Dwv7Ru42HTFQ
gs8EoqvRsx7wsXWF0Ywr/rC1D8fxS3deC92vYVzr9qWsJLIkhtSQYwKStiLYXC5lyCVje9Pm9bgk
neAZyOOGZcQhC1/qaouf8tR3KB3t41WleO08oV232IlzAdmO0TpHvOezjBD5aKPw/T7gfMvftLKp
bm+ytZlXrySkUwM/YdqQPBof+XdsxH4VJ2kkIkoNOTtpyU4Zs4gXXTkLuX+JrRahqcDRICVjTxOB
aYaCefSClS/oASqDiFJ7H8kZDE8otVjCIZ18HOSyZclN8rix65xFma/UIinqQkU59AyBQUIKFLQ4
Du0igotRhggpTQVV1OGJsFNM8FTVHstUfXgTkIRQ+WAtEkfROQ5kOGuNX08BE0C1YnUSilKKQ6aF
g/VQfB0HSvRMkqKUHW8uvmfaRP03wy5EVe2bZZTJA9GR1PfT32dyv7wB8APJssaqaz+EuxAA9pCR
XVt+y9Z/u0/f3Q1o/8tcC9f2bCBy8dSHasemIGGdWftA5TaZiboUSvgU5FJwlfWtbZoiEO3cPYMD
pBRCjMHpmhRh3oGI8Wfi7BMbfW6hf1sUzFpc7m/vhyqLsEvgRdKr6JCn4Y8syLrjUCa2vD3O3jVV
/7YItdi9z38UnJokcAFcHbOL+fqJKWyq44YSYBZ14nmStZ87RLKM9tneNSwNLsK5xfVDQAMHkMk4
WjXGB/h5VASmrE5xDsBG5UUwbiwhSMtJUQweoWHyhbPz1f0El8ZwBXBVp2sq+M9pW6OZ4zUaxwzn
kv/gTp/0+NVXuAI3GSRFpyL6ItT15iPUyYpxu0cpzu4c0ZWeUZppmxlcy7nM1RIP7swBP8B9xQfZ
iFBNueT7NzRHKfqWZzUGiLxmyPXOE5CqtRyPevh+21z9d70gF5/gHTsd0GLPoQZNE8/Z6+DaH+aB
5NdTOiUmP8T8uv41iXLp/nG0YE7EfvraqWxDVCMXQM4JDKFapC3+bEIlzpoPfGGZKSpPIlOtO6RX
2t2BUGNqOUSW7Lne3q01hqu7TxMzzpJDtPUkgQX7OfVvYiyrZ227k1Sc+9X7EhfZSEeLIIlqns0W
R0yFMN8wyJyahBkz1ZGaueh+oGZAqhx8rHveB1O3fgDy3BGNLHtWwWTKgCjMdbUzuLYcLLQp9IvS
yE0o5bhc8TpUmlejwlgdhsAcQxQM3nXtgVqNocl1EF/YTv4ouDsYLj4kRUrwQlJw8Ih0glO22huB
3lwnnEGsjT1jDPeGz56Veif/RyhQCXlnVCAuU0TmfIUMOyMNCciowVXbm4+7YSVwj0IqgkI9JpXt
91MP38iG9xhr1xxUXTEfMG4lmc6s4+n8/2E8sndrEQ6fGUNfphTPgkvbtSxpqRiZdtHusJo5MukG
Tw5bqSrVEke+OSkO3nybgUqOhdLMwsEEgqLB2Zp62yixS33bWyzxMniKOY71+ddxV2MkVLPE0kKw
osz7NX1YykmapajF/dyP7NnESb7oSxtSzt0TNVuEI6S1HSm20mVvU8PI1TdMB7DRDli+cKd/Eh59
ho2JzlqbwLyxvsxlnrtpdhNQWBqTUDpBCsCFUVIvoVStUBNKgM64SVcAmLnbee8QXpy3b6ir5kls
qTyCwVe+/morZ5Ed5Rnx4rqiLfeaNVYNsxzaPHNFLIpIHfIGJPhe8APFItW7VtYewAI8Eppel/jA
a/68bPYjVPhhh5Zl1ipuA7zJoVYcgeQ5FfQuh40lr2P9LknmYniQ3QIrMNkLaPUPxRfStOTp7Z8g
wjxIWpdOVFp+BgBPhJnar8TBXfj/3Jopte06Le7WGJeDPwIrS1h4T7UiVb/e280GmTe0Pj3CzHJ0
9uZErPKAKZiWgPfdzSSw8A3jDsNFZ40KKGIaZSTjJFnZ2GacNMa9TxT0qGMJq1Y7I68ahOJYWNbF
Y5+nUI8v0IIYr6HvpljZQeEExHqVnt+fpRbZBZfPULrEgZRkvkXh/4XiW+sjX8T5C3RGmmMmkIki
C7KDZG2p97Jj0HFoxrhBiQf99T/gPAKf6r/T78YRYl1/lQc3enlWMPJ5bKxru3XOGgp2MRr2qbwL
9gYVFW8ogKsIEQJiSDrdSWZJ4Szb4JnO5h4MvsrI0KJbKY7zf3qctk5tSB0tMzZLYcM1D4v6MuoK
yEX3Inx1ET4nq556xmk+dnOiVIZtUknMUSyVJ5vNoyvkGK9YqK6XgoATmKTRf9EtouKU/hqiwk6T
I1R9MWml7JWWa7zSOfVmgVCR0J/HFBLSmC1Uf8Nw1y/JmtCZZuZVP51cF28G47Jt0uV19BjfimK7
1YiruFDktIZMm1MuddRFWRbTx4j5ttVzh9+WPllfjdzuumhx2kvmttCK42bS4gAI/KDuPz4Z/kdw
NTvqhErydw+1TWsdHbnXvk77dQfg4owec+QJxtxJU14fmCOxXDzG1MYso7KH6cxybN6dFEMpL/xS
toBbo6hYp7Tbhwi8A1Q/e85Z7IIO7TK+BSYZC/gX+WyuIv2fPspwDwlSYb183tfUDV48JMKPgnWC
C2cC6TvEEvlqXxpsaKeL26SclLmVEeuWfIbW/PAdGdmlUpAy+aCtuX1AzNO59/tO2hNkX5FjOj5B
mxb+Q+Yn0Ml97KYVLzVCoFGpSp86ENO/eXyxHM/ssdf5YY8gbvmL5yLUZXAHF79+2+Og9jNMMI9n
PoLmaf12GH3q4b3cQY86B/n0J0Pdn80hhaSXeNpx+8jLpQlSCVVc9jhTejDc0VSYZljdi0LCv1NS
SgPr7GMrdQaJIwZ5DP1hr/4AwKML132JglAKfyb5+1v3tTIInxG75ZHK5js+FW86wB4dJ58oLh5M
xFdYEG7z7ULSLVSwRlj1po8U0sCx8Xf91oX4T60wDTPNimOPh9bBhKR+RTezu9ptEWbi+nOeg9Ft
qFnf70Txy92xZNqLKc96pfh2fFbaO2gN2UWYBy0Gj6QQkk6MBpgpyAEuKJtGJLAYK5GTd56fJ+Lm
pJKPHPQdfSYk1zgA59AmiRsw1hmWCb5ig0Ddl8grPb0HqgVD6k/P5uJeQjr+BwoucASwlCqnyVCL
3jnBzTgzMVVwbHH6D0zhIgnrip9epC2P3KwZ+e09l+wHKUmgiVke5i/T7XHkA1PnwstwHkxtRRaY
+Fe12Kx1KbbPM46SYskXrak6yCy3zm3A13LaQsj+ZIY2swECQSgYL8F3z7nDbVRp9etG0Ud6K0xv
eKuvTiyqml90SDl76CtLzfF09p6VrfwWS4CrdaWb5tq2cyxBhVD0LiF0m+XpleGmPWtmXITUp3py
oinp4N3R4HkEMR8phbq2MzbQ/7qw0D+Si4fajjwYBSXPxvJZ86mkfuVlvTB3t20VsYpql10cNjaN
tSiu5IynMLRSVtZmjj5H2Y8BA7Da+qIex4GZ2txpTZe0qNz7VXOxxoVumrUF3gPM9lJqUxrzxZSR
eElzm4NPayk9SXHAPhJQA1XvI+ZT6f6ruMa/Dl7mqoo3gPW3AJUxKrKtHuBzDogYocLv7NVuE+4T
xgFjUjJnotLNkbIfD1s9Cpjr1pmWx5DT0ntYojat0VhK4rEJ/+QlMWeIseSNsfFvR8t8RE7tKwLW
aGYaBUDOlVJvz1VJbMVNJbIwL05w3fq9Q3IDyazXbA94pHSl5jq8Y3jn+3Gq05ML7igrv7besu4L
20XkE2aWib4K4xdZUskeq0er7a2KommlY2ODnA+UC4SsyONb1VrfEEr/xLhOSCyfzjXVzkLMdxgV
Bhsy3Ze62mcgSAkaeANVvcsgWK+xXc+AKMAyrJsRsAADq2B/OgyRX7YcvWBuDxbFsS0GvO8ANowt
5RClHvZHx26LO2zib5YZ+kJK5uOIL1hqVjXVLn5YidYm7qjlOPTdwGkV/uw6qXJO99g5o2Abd4Sj
+EMIxCFQHZil+F6EBOvZUW5U12g+ZbpDCtPBV0el9/reDjVc5w1Oqcp4pcTy3dnLGaWg6I/ShvY7
apujMvZs55LW19u/T1BTz+5O06/VLUmN8ExpBg03ObX8kddeTuRFLz3laRwIkRl0/Q7Wkk7b7miN
Dj2q1I/2J6lbx20dvPRHqfzIWt/oMAhgwr6pwpkAUfV4NUApMlxvaaJDJ6ipYKpHU1nf5TfBGWkm
8BneFJgxzdEgi8BKA3ygUIEp8+3REKchATX3obCUSARuQ/3JUz3cc97NLVUfghI5VSCp2VeseBeX
u9GG+MQT6XBjuw9Bp8nH34QbQtNIt6ZRyygMY5j/vYZHkT5Tm3MOFCGN6vPYthOLEP3EivSvniTG
097imQ+pE4Wholkpnoxf5a8Jsvtw7oGXERRfmG6oGvhwhCLGqyus6C/k6mwYKwTaVB3WPqA393XN
fQhW1bFPlMKDq0SE8lJ+JUZ66JN0L1bEbbxOn13GOTtJJiuvGXO2rdr4TdR51d72rH2v2ddRohWF
NxXTxA4mHSuFwsvM0U1Ba6gn+IFRXw6FJsh5j7Zsh5WY1XPGtVgOyOsSsh3nH58jpIEMujs6qb+o
OYpg66rIv5hWYd6kKLl1FisDnivKOKTI3Gqg8jnZl90bhxCQvEWfF5GIiJM7pXZ4x6z0ktSnkymd
eBvUwG0ZXFlpTWV2zyUoe5oqnwgx5zlSwUiG14xNuJ9RrM59XjWDjZdAGaJdDpVTE+wrH3J/EKmA
wUCDpsUNFF66Q8SyNtkAJMn3rtkay9ETfUtFps5QopVdMeWorKQszJjI6yvynHP8wwtzpUeSUAHl
43OI11Qefu4ApaznSnnURGIeTEyZWa7EGLNv6LczvLQNfYVjZvG16GJgevK3AdipkYmEyt/Ws/fj
n97+TYbEy9cCxuSVfNjVyzFwUxr4cyKDp6SmCtR0qXEJwVepwFVaP2HwsXB4yE+prQBldjZGYe/9
yUX+yqEHB5Dj5zlBQEYx/Y4DsZUr+piKRpm6Xfx6b3+vVjxt7UULhJk/F2p5ghT1JxsbBxqRsX6v
n3Efts9E2+NccQOXnbaz3GTc7ar7lH9LJMSSSUtnv2yX3hSPhVp4M0y2zaA9E3RtF9hC3D1sH6d6
2M+8WKZaCuRN2gjHfbQ/qOxNsNjxma+0rXO/EYOFNYAaHk4y5sy476c5bVuEGKrNSUQq7xkqQFdl
Kk33zhtmETg41j/ORCB8aVwIhlmlsoNRUWS8b6qZcgOhS78aPj6scUvgqYSruqAcT1mwSKYQHyZy
FrKWgTLX2t9ozsZrVy8ldGTaFsRX9cDTQ1aLUi+PO9jafPTWZ0wKAkG2M8iGue1xRKhy8dVSh5sf
6Lzr8dAtakepjU0+U7PaRestl5KaKIxOo2Jz8+bo5b/lIBnG/Trz+hKHUm1siXELs/M482rRZsW4
9cTdkt0qj8MdTAyrH+RStKMGcwKsml6r+Bwj4FvmLDqbusjNE1I67QRh7qpLFR4W3qpMYSgaKz0J
2tKsEwSswRMzRTBY1Iv1URa99oaizk1JnB5AqWkp3IaPu15dcj/0+ADIjTOFs0MzTws8R2r4k4zh
1EGzcpI7zwdNxDLdVfBTlNh3CHW8J339xsZiSHEsfxiso9ConE7T/R17i6DuY8uOuDOUIO/WFklC
VyV9MUqn2mysGUIZkXcSHZDx8pO8Y/jWCx7oJQTVSpEOMyPI1Oe0qk0vgIbA8IUKGYa9kkst67z2
9Orucp2rFzjw+sMR6SOYsZm9+ban7NbvO2I57nnw7JnIIHfvACQgKN8ST0slOqKVVtb/Dfb7+xNp
dZkaF717szTD1RoIfsqwq4rflv7Wmx3R2oe681nD7XQpxhHJ+EeisEkhhmdbAYuztT2P3EldlpuX
wW4RtXkV27E8qjRZbcyIIba8DgpFENVEbnH3PBwV39eTwZaUdNuW0OxT2wNmnlGpmlKeeTpvD1WL
jr3pncB/CxMhqQLRjHSpgoGr11VY869L4xHBO2UBUif07SR4iv85fpr0DHdB8qG+YISM1OnaTWp2
ByFEuZZSPCktcaOB4E8ut+hEUtiUW0C30bf3NUEyG6BSSeaKhdNYBc2IH/QZFmFvvbJ5lY0ZRhsI
pOZquTEAAjMxMJsJLBCInPh1FzY6JandiMDFSPEHERBhS8XdPPfw82/ADaZhZpXp3tMvOvDti15u
9ebQFPDisdulH8gIL3VkXRcU3W9e+LT6vPxvxxelxdZVAHeKbMXwseMxLct9thP6VG8PFDT8SV+i
yLXEEM7lfw0lX4+Q4AWEt4tYrQDY8FB+FKH/xXWfC5+soMk0QxedWVCzAyRH1SWbNAPoRsm4H4n5
z0hVADdVmDFco/bchQPcVHNBvBvVB3J1AAFvs2ZG3nCdV8tFB4Ygf/6bHpJ4gWzmza9ILmX7kk9o
F+fF3tgNmFviujk/8zSbo6O1i36SlaNhQVPPZny+mWQDw2iLoFA3c7SkSe02yX0jTLeOZfGR7JQd
NpYNVnHyOGYlaWehzDhlOzTDSN/UqHXNedWG8kiP64fnLGA33tXNrLyUwulbN+z0LsHg5YyYUAAb
oLxtRLybU+buwp9C/Y1XS229AES1wNNbOvp+hADHTRo2WBGULX8laA/YdBErBX88Fn2pPy9zU8NB
dTMaG2azAImsSbOgQ6kUvPx4LC1/6v3MDccTI2lGFZfqRa+6M+BG8pKssqJ47lzqGiaDyegD6Dmj
a9ZY+wLD4CWwke7Vis69zbXA2Iq+1T5/KajFGxW5PiUO8aHYHzlpp+cGhWfgJJYYGxxR3E41aCWD
rOnZ2GbbsRNXG+NZC+d49AysU0U75c3tn9P5bqnH9hqI3iW6eOWNKSJvWVuKPkwwD+UhZ8sAjGE/
MOCGUuY8x84FIqUpXWD0kc/UnwEg5F1OEkgiBkG02/npwAlyDHkv+zZ2ekBR3FLcrluzh4YgmmmM
meO3VmF+jQ3CIYLvca6OFV8M0Yy5zR6FrbcWg0aT6M6sZaEOXmAuEZEH9FyosaSecbC32teZG3bD
Dg3WvCDjmMyIjpw4tc943hzKUOImfLauFpBF5+JczxHzB8wOVQdmKE4LHctm/wOfUOyCAWdDFsWx
UqF6GjmcKvFsIe+IW/3q6Zc4coiuoX+dowKBt3SVxF+XWC+Oo4qVK9FrvhnVnTR3P2j6tS927VG+
DIHcaESHSIXYh7qDDHuW/Bxme+c4vx6e9qpWqtxhJ2a7koKCZrL+6tzeQxr8T18kA0kB5cofrxin
ntBGwhk88yEHrDP7gcASyRNa9LPPhxxaspX3HqYU7aWGa4V1e8PtDDairVN4fqHkFjWixOpn1hv9
67+HE89q+mpsXM+Kx77qkuqJzAtonOmhokqPRUGoP5vhDiahzaqfEt3b8dtazZkEoLs92y76FoO0
GlkOGFmoC//9fhtA+tqYsexAV3czDPHI5Q/39ThG7v7TUdftgFZbc8hFbtwtYVrP+i3HL1w7DK9B
A5VNki1xzPydUqMRf4qj+0fi6CPijlVHZY0ggQMgR+ihCA1mKa3DqtgCTVjtek4JnyHqL2nBkxfq
qT+q1jYlhjYo+C0jgh4cXAFzzjxklT4TqEYU1YAF4VnkoaVUrmbrdM2n3/imdxq8lUjrDX1T/yJA
Po0Qj7xhoQ7fSzRxAkSCuo1MS7dSdp4zlx1YKoOiA5x3eIxcqdl02VggJP2c1BAm3JC6sHVvKBbi
9cbQ4wYyHHDtcwuBpNsHDEmqRh2lqWL1+f/IV8bZOz1wOYVSo6ANAkFR2Nqb1uaVZAJU4WbmiF/7
g4zkgny2Ahrw3XIYghXCVydapFRSkNNkjCMZID9hgBy7P1UcXHre8UbSuRa9Vcw0Ayg7IbqgORs/
6HVABbgKjtoGuz1R1XCOEjYygGNjBXLI/c6eo28HCklEDtX9hmyUNt3RCk/rVSpXn+tyrbevjoZ2
ORF6sPXgQJ9cFmEx/EJP7CHgWQmbf2h7dLWzx3XrfV9Kr/IlugxjVqxVDfTcJm7d+2WqlaH3OE62
O5C+yoSG+WtWKDSda1a7ykuULpewtuDUTTg28LaHZdP13kaevywRkyNU1bnp4V1htLW4LqZx7fTq
Innx/++52lqZtbwjAv33N3WGz8js2xHTOhwaKDJ1oZH5b3uU3Gf/KNk3OpK1ROe7ApKt1sVlDEjW
7oVvtD2riTT0/IfAABOzRrpzyZi3wn0HAoH2edu8Pvmq/Iqyzmhqaofoi+1jCjQnvhuHKmc+Tokd
zdh4JN+jduUv+meNAiwlUfFbG2385BjErgphBrZ19irPjk0VLDo2VIwYlrJ0x7MT2xWRKdkXAEDj
F7Yfeo4btYLdaT3GqsznZPOzN5yG/nBaEQJZnz+CTqxJLYaRUZDGOoh7A6k6Zz5BoC83GyMNJlTh
d7nFMkw4QuT8rksFQsDTYRDe8hn37aakzZ1nW2hrVyPxh4oZ1ZSqY2DXj4eyhSgS8TpTQIZ242e5
yEendv9HM2OpyoFLyySAe4uXawIka3xwLBnR6mlcZvQEyHtAOBuzAQ2/SImobz6gg/o+BrcXBaFO
frbb6ZUubecTUkresSo7BQCxdI32JOoUer6PPws3CNLrUP9HgjlsUPftBiC0Rm/v+wn95TnVzux7
GKbA2k0uNXqzpKxHWTItuuR9NpHuT+pL7DT2x2fJj2ca2u20bxWLjJLF4gT3LVeUqQm/hl2bqsVt
CinO6icRyTRXA82ZE/zFefqESLT/X67NTtFiwClA1dCgRT2/bPqrdkLUGOdLsMPtak3uMuTDaNZQ
NeN6xt2cHaYefHj2LXzUyKfoHf/Ota5DnsQC0xqcCvEbr5G1PznVifxwSDbXstWNk2gKqbPG8n/b
bKMcRBJixH29cAR6rSF0iraBfZzY6RxXJPo7w6cNyzBCnIPBDCDl7yjFjWlaTmVhQp2aaIN5IAsg
UqRhOPipwn/vinEDRj02w9r7I9/wB8+FywIAjP/fPLgrw0fkLnLAEw7JTjHjS+ugIAdVZSG4eb4W
JB3TUCNIiI4qrGrk2FiedDRk3kH2NtJvp+zcN5AJpPTowIuJo/oWCVqpbCSk9pD56hr6xjVL6in7
3EnWn0+PpreVWSDYx76G6vJIk3COKqTGwijrwEyhl46v6YZTXqEf/HT10092X4IKEtAf3iIToGaQ
Lz0bbhJ35Kdbfd9q8wBC+bymNKN46bcicW5rm9rGF724iWNjaoZfYrDavieOTAz46HP9LAZLzZXD
ABkvkb1RAsUVnp1brSDeJAv6YM4sdMM3EXLyfWlM+Axkzpl2TilhYL8Lz2uOq5NhibUnNTeVVu4K
L/DyJ6tVcSDR+DZMD4dowdUIVtk+cobt4xIguRVEuvppLXGG2EhjRS8IqR6f53jRYBAFsXoozI8K
kp+sW7zPZ0+BI86jk3wNNpdmw9g1k8oUQZvNoe6t82aeLz2j+a1lNXldaeXsYi1hyCyKqp2GqUof
OuHvNAibK0tW1nosmGaUj1MS4qy/igdFEbsnBcmp2aF/s78kb3vb8l+YVHQjoA/bMENeFmJ29hdN
1eRjiXTvUMAscDCuBQtw7T+F6AcLI14OSpUrsSKei8g8lUD+r3ouujaQ2lvkASqHGc0+HAfr7IKm
gxB85qHi3udFF+mtfL9DerJnJFGTyL4lLmKEr3hccVtVWtHuxqmyipjpmTKAEYAL+XjANPAvlCZC
ny+Iuxy3v/0UmcJLN9nN1zDP7J+EkGR+UdkGFlMRZmyL+J7R61UAIb9tws3Eo7bPycNgkIBxO0Tu
acL0ukS2m6L83Bx4Flsg7dVWKzmS7GfE8HaaAwBgMmA42WqK2JT0ySxmC4ptR0s8aq7Xq0nf2wzI
j4UhZ9pGw6N4p/RBcEuKKyNx+feRnIAHMq8g6D6zOBcY3Zs7k/eGdOFLcIBLi43ohHkznrXFRSoy
fBd12FQQz7MVpci8qiHFDgT0kHLyraTj+GzuBwiXx7jJhjITBFAmi0Jo8OkUCY9L4WuNlZ7Q3bM9
12LU1SbbWxZZS3l6GTiFxl3I5fWUB+y28SaQjeTBAnZO5naS2KZ6opW6XPAUErPO+0WVa/yC3Lh1
VmXKxAMyQPtf5uZ9ccTj4sNV16KB9OeDLOaOPORntXrch9eB0yyMmtrPhlR08WvMyT7FSvQwPlP/
qniv0dkywmM4BliEsbncPOJ7d9iKTejn2Kl1BsJIurBgmXy23jOiEzTEVz9ZThoZXq7zcBHcfkU4
e+Fy2dCJUvACT+x/FYDSZdQq3epuHs4/B3YOf1ZYFr2HcoYiRxLT9IWz8JoK0LXBHvpCQuy3nrBy
TYlmW40EDpb+qq9UscPgnUakrt/2JPlmsfitkQwLWltpNFPJCG8nZ2t5kTcxJK7HWkPkOxUD1rKf
ousxA9tXyP0BKQETp13U1Gg80siBOTC2QxU/fIfbq6PCx1KHpYvRlhiivxhJACU8iPx5ktXzHOBq
CABbLspkF01HNHzcuk3lkzl6ebnpaLPBRYTv/mD/PmGbw8mMX+RQSJ1vx3PkO9Th7Gp/fQtR2ihU
7NmPhaLpi2hvH8V9RFd97nQFiNT6QZ/JcHfwwA0u9rsDhQckPNX0P2XXblCHqu/Cwdgh2nWaQqjt
mu2+CkU8nWro7VkoDR26lyp+pqevCkS0S9phdXlYrfd7Z23xJhJKAzgXzO9lysqJTh7zG8aZbvF6
D4lZW0jt9BoltiBrMs7udcIhpYe01cSbdIGzS8alzvqEIklljC6fZqZOlFGcqwuRrIZJhTQ/94M8
JmfUW4kERU0s1yWAcrjTHKxM+7eFTQ1upuwyv7FF7rJ5HsvaSx8c46T0dNziVswFExGC4Mec2LEC
t5RSjMpHKJyob5/06DzQR9Z0KPmtLL+vug+HNEwCD85MMzLS/9/SxqyTj79x9n7z96CVsKJukZJd
1QLEzLAMHupcSSgAkLXhwXH3phSSttPY1B3t9TSolX2i1lq8FbYTEb+bKuSyp46yUV0V6g5FJ880
kO07lTyQ+6hMFbHNbOb45scB7Nm7cn2s657XzsT6JYNgI8vCMzSqF8Ys0B2SJWMj3pblyjaZN3f3
TOyktLe9UB9F2fAiYHd7kJHPnZpTB4FGKlBH4zaYo8WOhD+E54zss9qhHvCY7x2Q9TpYNN0jpjkJ
6IOeIlplPYFw2mk79WTKihLUiWKFA4BuFZMUe4Ir/P6v1QlfcGGuOKEIKfTWc0r77tui9fDMBsEz
ibYxaOrr/dLT5bP0h4kcCN3rdeoeEEbN1P11fJT/v93jFeWLWMYiYtnK40tyyFPL1N7j5XVMLODh
0J8+BEyaTX3808Cz6zpziaOxdbI1GBs47A9Lw39QtTEXyFyE2MAfDCrnp2XwEYZRdDghavX3Xelv
170Ouw9zznsqZwHtVvS2pd1PFnwFK00gKwL7KUndL4KA2HmII7FA+2xYL70YemeRCBzsg5GOo/GV
4wgPM3CnwPRyVtTu1dEGoEDZaGh+bhUt3xtJgEn7KikED11+Dw0YeFlSunE/8vFNnNpA2/WYUr4Z
Syz+Cf2tpAxberICMET4zgJluvcPI3BTTARP/80oiIK2EdrBtFxwQJKuufrRQvNnJ+UCoTYjWKRw
b7rthR/RFHsaYqy0fx6ML/GTC+9Qmk+oURkySs5iVKyu/LUh7jg67CR+owwQCjjg350F3YTyYu6l
CT2n8aAsu4GI0dSR+ACoXpiBFEuQmyATqG+gBejCcyk4t8sU/a/gXlyoh1xY/3PUdRXGTpusIiKr
K60zeCFwQ2I5wBg8Tkh9xFeLSQfUreu8t6d+UDkWnXTkZJxyC7Dz7XD/BuFDv9xwxgHMumCcRJzq
flYSud3SsQQWITT9qclvyb9mKQu/BZfZw91zUe259KqXOVLLHORw9kkB8pVqSCbU0Opbh8L1hyi5
INBx8UT04Ot3QQH19Cf9OKT7UoWDgp9000BMv3PjTJVHvC6bRH8dUSa5JmEILmHsc6r+VtfvOOej
e6oSXDKBtIOXCbMq//cEJRkAuUq1b+Ge/gIuA5CDrmCspDngCLaIBwdxf2yk1oKd/WdcslCZJhQn
x1VvtGnhontDYKOdYJGAuGVmAYLYR5tNPKWsuxCM/KgC7a8zFe5SJikjCYP227JxDlVw8b1d4UH0
7DpcD05P6XOgKE1Gr81iiqocpUWHIbWuCSAdJt/GApUumnbch08d1hZKi+LrN+L2Ihwu/fDp9jNM
6VHQ8yS2h0tPvawYDmhsK4dvG3/bjzQCxDfixrb5iy/aglPLNvVukfAMbx1Bd/EY3AwNec0QiYYQ
ZVHA4IfRZBTyTysAOchrRpL/XPiviVg7whuE6TRfzN0XpZc3gJ5lCyRwwd03oFt9TUFSkebcrA8M
MCLAFYHhaOz9H42jgrhnPCH5JmiCJgqP3O/yvrkuTxwwnCmzloNPPfKZqtiN5q8Dwl9i6mQWcvGp
DEO5xTCEGXRoDDGp1yX4StjqK0BuKYK86ZOPh7lqPToWVI/kn3QFFtjyk4xGb3Kmfq2UoaTY1+EE
7h/DVUZahRoZUipw6i+3Lbt8EqrzUQT9hwvel8mi25AnW0ciyRL9/eUN1297IvXZmZWlK8fBSIGL
moUBdF87j7salcBxrWpR1Ao7GYFvRmwWMuusVYCpuypm44oKYfoUyMANwHv2ZLdi4gSdUp5D+e73
0UYixIOuvFTZsHhcb25CUvmYAfcmQT4zb6ywjVPdB8KkaW+b5buooAPOrnxZde8Ms8c4g3rRuw1/
8iVoCQ/qpnYv1/bauZbtfSn2NYPWIi71Dz78HAoM8QpuwcSNTd9Wy8DnvT+GxYI0p1BEPoBVFWiK
3s6jArVoKFZD2/AmkjhP9OePuvDLDfK/MmIFfKVF3i2sUlNOiyFEcFjHaKOrMsojXuD89IYhTsoU
CbSXXFzzxcU8aWlgTd2gXE3+uh3n3fmqJV4pZT5dI4kEdbiCo1riIAJ1mosgi18j34beRC5zU7o6
rUgGkatdnHOKztFeZFApG68/vjKdM0HEY2sYAQHHT9rk1M8qSBjKCnNwEd+/xJ/L4/F06kL7drnc
/y/Ty+zfzn2k5Fp5oZk0+lzIq+UrGjBPAh7coV013eQuL9HzRQqNNMEYfhwYw1aYfqfs1o2W5NQO
6iK4mUKYwQY4IB7fYZ2+OBxQ0NewhlsgDCAwUC9yOLZQZGG0NJvo4ek08F3CqKjA4RRoMicFnBKh
OZtxmVcfugstDhUux1kICqQp/eKwBb0c1vH/BtOoMeTIPda8PmTjRYbsrUarMunJ3O9qVcLPaAmy
w4rU5ZWZy9D8Z33poDrK3cD2qfwyHs9/e579p4lQn4FEYcyHya7m+5F/p5hjNuiSIh8jsw3jwMN4
zhuze7SarJplX48X0E0YkKZ2AHf0iofNWPXO06rmo4Rrgw+DTLSnui3E1ERPOyALEr+NqYVONent
Dp7AapHM3gkAUk3yV4TCZZNmUDuQBTLGEq9HbX3Ezn+Z0J/gett8s9gmukkTatbZYmYwyBI9tOie
v9/zyMI2vX+xyES2/MmdNDAkFKoka2Jo6VJAu2ezWhC//uHhjG4o2g82UB2qnyUREmmH/6ExbQH3
pEengHeESlA43c+uiPAnahG5DkcjucvHXgnbTj2Hy1J6lGJhGlsh8D8X/1dbRxp6yB2VUvdHCnt8
D/rG0nnGzFHCdwUNeKgFJ9tWUC5ELDHCE1EzX70SypBRbvgxUs62n4bXOrx6TEZmz1r72XS54gAl
lfIuB+rYv9B/F6d0/9RGcvIcSWZ4R3niqpevPEKqsezkp7B7AGYzcI0zxuiU3pU0neg+OwMOTOxA
G0dHwFT/Fr3MjQUJnXPUC0kXFoJiaLT9FOhHzfr1COwqoMc2rqnbLbP7wRUh7Hz+Qly432ZCZL0Y
kr4D//M/eISPe8IOdp1v0imYQMpdYBH5d8qJeGW4QgYTJR4bCggAALmMJ4iOiCPIGoNxoBydYWn3
TjK8cOCn9J7xZw/uBapg6ZDsMnuA17CrRLNwIKOM0u2wNd+KsJ5ahO2rlYxAWf7grjUmSbwsEMpC
0VkmIY3xAqbXVRHBMbGdoajf+FDim7LS3uyedkmk/XhW2JRTIVm442FAeQmqvl+MRV9NEEzhFE9Z
HUvBdCTkX0f7FhIGNM5PL4bKD7Vz55HubcQhzDj6AQyGt1k1j/bgdlFOoqc0evrLbnqIc9ORaljB
9jFYrfG6heAjO+mIxf4hWc97FGv51441XnA/8Klyvn6sK7s+/eTyYvj8vVPTb3Lr50ZGbXg+Xr7o
y3e0kFKvN/QVVgEtBjXtNGq8cyrXYGG50phkeZtXK2pEUUzzvWLoWnZL3fy3kLHI8p1XOgBUDJvx
M5Z8fULIrJ8PEMEiJU7nj2/buI4fkKKvici09AIEcyeTjBm1w1nadUPETt1htCJyMilYWamxckUG
xSZ05zSWxbY9JGTgB0ti+8SRGFaCijhBeS/dtNWVjdSQYfkggCLoM5FOsI76iq9oEj4cOyzxvvTq
Kr2iA3ejqeoBvUn04gfXHavPk9YiPi+QfIEyTQDYH5XqBnf/k29ACzntV+k96Lv2UC8p2I90kII3
PsMKY14UqpbliYssmQEICwphi/NNkwjoNJHFtE3vQYWg4efY2FrNG6khtjUXFa5641I/RGaJE2Nq
2Zo36UvgwhSwYf5olPAs8SW1gVrJUZuapnZPd3HbfEOcZeJJnAhRzzwjyTrQX43cMR6w+Ku8eFr7
DQU1OpsrhcdclzIgXjEBhvMaHFI9LpKj579ycEwL3Nz202BFy+495zXVBhJmquooKuTPHSmdJhOO
BaK/qzF/lM/RIrCbuFVR17qHwkzE1h32+cBfj1ssujFT0aacgx1vtaKZbaXzCIIn6pVO/V3nSrjp
CwoVNxp5bLT1Usokbv61zIhGeLAAhpnur5hvxiRR9f8fFxpe93TLF97hYe94iUwlvI+/g2QYpJSY
LOJTpr3P8nNbzKFk2f1whPBVX1tqVRjQ+D8Ax4TdTSmSxiimdT6tOrYebEfuaT8tSum8cvS+0M+8
4l1QVBTH4D1U8ADceDEk3UlclUUGvhtcLqj3ZczJnjQDcrQdJie48EF0s8Ea9Asn7huI3Eytb5Cy
AgEG50EJPy2gukJaMgQr6UiitHxx4a0YRVlNWWAP++NBniwvE1oZ7jYWihZuhkLn64wybQiAk2dS
vkDOwbpFb7HMMq37eb1iAaBQYPpcTqnetwEalv80657c9w4XXREuFBus/mp3tynyPphEkx/e5NbC
Y6pohEZNPNuFN/pT9W0UR2Iwvd+D2JpUGnzbmuuCA+sHp3vT/foQGhAuJI2713mGYT9wHbd4RGmo
Lbmt5VZiHsh63m4xckff5hY+IfTZCHXT+WVadry17awWIkeo6qGRAiKVBbFwLUSuSjKPrx0byAii
hsV5jcvjBO0UXGJvUqdruaY3oA2bkrDzkUqJw7rNT+gYsCQuDZokU3FngH7VpH59yKYKmh1eFkWz
XYAtoDH9sBYA4iyz9Z8XXMhrWVm0KDCSqf3JLVSVgs0brzz8aTwwyFU4Jrlg6YI8M72GPAJ/41PV
+71zPPJtptz5bLjoQeyjefMDRc+i69uZAk9ubYeokTfVMDyQuTAl4BGAZktijB6iIlyKvGfw65d3
pEETZ8ljYCIWXJjG6iPtKclRTs+AKouq8jVW+EJwC4qCWc8Wp/2hBsmFl62YlpUfqgITFF+f/zJi
iTW21ML2nMr4psZWVXKIgx0K2WoR5Ns8X9mc5GShFd9Z8dwHhJ5be3xrEnIwJmCxpgyAugohxFCc
H2WWrKMQ5naJM6lyf9CnDveP7rLKWBzXbGXyPeNr36xAlgq2SWNM4WcbL4agUJqoN64m7ukUr5jh
cJyKKdJ0CZHWNOJYvZJZwTHlGljFBdXt1TCXo8+E9NC/Lel02yikvnZC3/ODmymZq65dncboPIIk
iLW5D766y60y00PvU4ofV8qByndHvTu5/qpBCUgdgDPLIoG2GBjODumLxUFpHeAw79rRv63LZWcp
aNOyDcBe1u9z4SdUXrcTrtoIzV50Fqjb2D0yHd3YmFAdzRlcS1q8ZLoTJd4wXC5N3ggBGMeX8EZ3
nRs14a7W5K0saWqiQFC1tuA0g2NIo4Kc1XzFEqNfBtaut51JiPfwMHJ4Dm/TCTXZAe2WwNmtNstQ
1R7LtHNuPx2CxU2FMovQzAELgb1+vyT0g0kuGUqxz7BKTq13wibrRobjfFExKAJQICVL1BLcDu7R
9g2fyXLSbUx6Xo9f/0detbA596otF9vynkTGE2EESFfKZTr5uVzuB6Efo6PGD6wugrqSOOMoWjzL
AzcMAjCEINRlIspNCAAFxlq9NKjt6pBfTPj7gu7xiPJZ0Xj6FVhNSDdk+hi7OjA/AcvY48lXYq6l
2gpyxDOJ4OvuHll/sGMOf2cjJ4DqgLxs4IE4WLNLCAVWUYBwzVNkq1kykRzchZj+7Q6W8eYiwP6W
wCY92IKFvRVV0qoY9kmjl9QTfKM2h8rACahFWvBZzrGxs2RMJ/57xjMak5dmP/n9Rn7ylMEFgDqD
Szu0Yb6f15Lo7eUIsJHUNaiZisHIyQYs41ViXDXyfHq5oHRRs3lLkbBdTVeXXrQZIgvmpuv4NPCQ
BZsV5Gr6/BLuklVZ3dTVoQc94G077JnUtexsoHA/qzNm8sAhSQkeiT1DgX8FtpmF0T/vZmIrx7gS
VgZpG5i7kmcYBxF9vqz6oJ3MMyNxdviuCoCPiX1UrQE9nBFGhjWbAOgLG5gB7UV7Tl8An0p+WFD1
dXrF7MnpAZsZubW5km4vO7+OD1gnlRNwXl0GZqrtH01aVOjMyAM66vIzFez5zwvGE2BwgCJNuBcM
5op4qCGoegDNEK+WfcRkGY+sBii4uTBgmwxjsr6GfvRyK/FBiN5E0gsbXjTk8mBONaUaOjuNMc71
xL8r6tT0xC3K6J29lF2Vlb8bBGtKklhLaQs2Q+7Naig4hvG0ZG0m0Y1TS6mpcxew/GzFm3F2o5m2
98J3Q1i7BiiaXenGGqm1nyh7wsEKs1DCemLUgCht1VPUSyYuHma7mSWhbdR2Qn+C3P/4Mm36188m
nyDrnC6ZFWFB5EI/CpYxFNFakTpGS/FVAB9PDUYdhUvfz127honjiAtq5nwMPEI9WA==
`pragma protect end_protected
