// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
D1UC6C41p33f4s4GoZaHnjOz+AkRpLQuDx0V56+18sAIfBrzYHWTow3adpp7c2GsUTvkftpXCiYZ
cCI2co1bqiFfUgw0lG06HBX15wLdDDiAUnq1xOwUbQ+eIBzQQug8R65B/akP42+tR3yaS1SdignE
lqdlKYagv4s4dP09FcqScpBMCS0flDmQ+muicxjQjBR1ULQBLnQiWg4YoakfXMvm5I+TgTU/TtlN
tQ9XS6P6nNv016uChna1jW8i65TitHLlqIp2jx7gBHpdRedab3nz2MJ8zjlt8WKa4rCp084E4GFW
6MiT1FKlnCNF5vLnlzk98DeTTcs5ITjgWg+LWA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
DJ7PF70T7K+NK2ThVL8F4awXFUIZEmi8YWXkW3gyIbhe6uG4Gza9yaaEpStSrfTtuib/nmcU/znL
h/i2FIm9zEf9B25MUDg4989tf/zL+QZvtkEWs/52Wwqi8CRMFWOrDF8uEqS8db5YnE8Z57UQSfPx
oQFDrGgFicR2jvZbY5aLau0ClC26vf9dmtLQctSwwOWCVW9xujNmnFtvAKZ+/wqCU/d/mnpOvjcR
dMu6LxqyuyyUCbTOCtGnAmuXyo1UJsi0GINs8c6cbkEeNvg0BcClyysNQbv5votGb/PHbKcqwtfj
1FxjmqPITkKenqKodZR6gvj7QUGHsYwCIEwMsJzQIgZuhVJ9X+yLAyHYDB8W4FLKgN5vY4RBi+ld
oXBgO9OR6ExtcLMH1G+og1ECxR+TYcI6zKkiUYGWkoKjuMNyUjdQPfWnDKaRvIXTzhif6bcbf2o0
szqBl1nQ2S1tysfsIMcwFFDWNt9X9YDse0cK44B5wlZ3aKMA8lSiewBfDyoY/mWWvOVmEo02ap0P
IS9i7FJ2jxnVuRHFNISmjCPCwTkpE++fwT3XX57lWA8fTKuCjJbhCnN72JPx7/ZP5PeTbnNZEBvO
6lOTJCn1t0/j9NBG2Yx3vTCV4wbX62Mo7FgeGy8UTh8sZ656XFI05Ilg6u+NeKQrAj0SOdHy/7DS
SVtkNwKmtF3A+Dcr6302+zcq/3/ynch0z1Cbr11OHlcK7Y6T7AOjRYgcNyI72Ph+hA8dYeOOqrgE
d5TJYAAYIZT+zm1/HW1fcRl9qmrLaJ50PV/xmqI4LAxAgMuvZ6zje9zgZIr2rMHqn8ND6HxWRfb/
XL3NPoAa5zvoy/wPu1h9iF2sn53zmSWE63dHXLl7Rnzo/uTf2DRQ0LzKvSJCAYEa6myiLunZ0yYv
djrBH3OZMza/cNdUlsr4hCFZATYYrCVqmOKuWOSV7bd9UaFWn7LGhan6c5YZUhzTQKkaoOaXU4S9
VqiCh5BBsRbL/gAIqL5H/crnk4w4io2iSoBb6EnzVeN+KoKbZuxEttSDAjU6Ewp8G72EmkeW752x
X6ZVFPPawiCTF21mbhOPN5laJeRPFH7HAEKEfMLvf68X+hkMHXNxUg7Z8dDNVbQ2dP/EIoFcVPR9
6vujs8QvOi5AWecXQ67LygG2R2g0vT8fZ+0jlSg/WRbfjklIr35pVqxpDRAKxdGde+qrD0IEk67s
GAQh4QxMMRnPU6m6iJXdAXg5vJZNgtVkdmsT+/SPvErirp+1KFDYWC47TUdhtktfQLXKNOHLtQZR
QsZaqUGv7WZeDirXFYp0Gsdq9vuI30QCD9fZaFDhz1O8wSpwe6NV/K7lMazxaXe0M/9f1Cz8ROcY
44B9ETCRoRYOpIoyOFrLaZkuNVVHkooyTVCNjy+vcZeKs90h4QcKBOfiLSMpLx7aFsYsu4DhdTw6
8W034zhwe9IDVrIgegOCHJ7YFHfuCBrrIoylMKlzKloJjhBkxy0ORuuWkC8d77SfRSZa5Y1p9L9n
Aok9icEhrmccAxY1V83ZuMzWrcxMhUvjtrhyOAldqH8068uotjjVbuehp9/7fqOtASxSuJ4RO+0U
P8XrhvlmPHMNtYIYRhM4opKsar06GEmqlf59kiY0ZujxtSQyIUKYDAQXk46GVYGxV+3Zp9B3X6Ny
sjI4Qyggq86j66aqax5c1nXGwfBB0R2VzOG1Y9MNFOT7LIjs2aHSXOW97tXadt9DwshSNPPIbgoC
BGgOx9aX6G0fpS06Y7LsW7pqf5kDyMEUPVTV2EfkfRLll7xcOe1rDAAZhXLaY5enSNIMhmqTSpOn
pKhWXJqACWwT9ygPm/powkGv13IEWfNEuSzVSQPVbmbUFVu65SZPKsRqVCDk2pUQ1By6gccqNad+
+yHdFFtk02+W85GmKW7JiyJvisNoSwZ0EVmQXrPjsfUpvFeNM2EOZ3R6VYy/6CjkQthSHxNqlOBs
/tFCkOm+YoKK6QaKdrlSepxywZurzGyE3niZ7z+/G+QzeFhSmOGgcWIafSq+tbrzNivQqm5TUkBG
yJrotnyEVJOTnwgsqRYyc9Lv5itK8+gNG5dZRQ/tWQ2YxL6r1+qOL3QuUjyXPveebD7tlxko5ecT
E2k2ud1DndCtDeGFyc+4JaPaN6JCPUpXDWLrfQmc/LcaRiatNOSYzlYeRag65yMVOjTQjL7A3fR5
xCs7Kb0mGEQZPJVCfutiL66il+37b+W7r/jqNQctTAOZZ+85tqZ13aAVq790eZ32J+7Vqeu/9jM1
QO095IzPsaj9ViSiStkxVetP/3Bw4EKW0jplTGyKNE6CEoPOg+CGgJzQgguc3VC722vmm+8fTpdf
qiNbbEkout3OTZf1ECKbPooH9ihsxmg79lSykpxP1aZ+TzZ8t5V1j0Hs1ioKF7BvXVKOVY3Jj5ye
R1ECue/hNfQHUBu9IHO7au5R1GraXE2oZGt1eaYo0rmuLuo2HPc74skFnDXtbnKSQGMbq6BZqU1e
6ycKYTCsxDEWG7VP2skJOvY8W08NIYbZL2mAGRc1aI73rYhvXzDyiswDa/jdbY1rco9rm4vVTzTj
nnaddAGjxX/rQUEsCT5EDJ6NQ5KXGSdv20prz2JjexISvybRZPzNp8pn7rRUdiXPXymQx7/zJHZT
GPvv8ujY9cDfcEwRVunj0sGahkYRGxZlzn4dtKGMdr9iU9GyUM4zEFyBdksXMcs6p+opnhcnrgpx
4aUEAR8Jsz5BnpG6hu62rapFF9qyuUJXryAn2F1J87ItAEv+Jk/rkgC1vyaJI3F08Fi3U7cDMyEc
61rUanDpeM+OdLOPTOloPTX9kRETYvmxnI+2Hd0vTfQM8Zmg3l50NPQZMgGZei4ML/qIqa7lYktP
kfv/uWiOPKLlAerAV3sCZUO7V5Flsioav/bxFWySbqn9qQ5vjs37Y/edrfvdhHLV3oltW1L/P43j
VtSwcaQ/D9ka4XsPasEh8terX8fESgj29A7DCrX/LUGRspTa0nVrOjksS2jjdCRsZm09hmh3nqe/
nfYeRjY5gDM4JTUA97RXTXS046Pe1Jh98mThLEVsS8FBim94cBI80TCsy8+aLLa5YrA1LOMAzC2s
W9VyUN8GHBgUguEthUzEcL+eJJGdyHlHUpHagvdbHSJMIzoM4P+IWc1EXUigc+VAtcaS3/7mYNX0
7Cy9OjLBav1z+dITEedKhioparvR5j9aDX/oQnAjTHWEmrb2DWLOvr95HhTU/DV3bh5rs+OpD70Y
lR/PAKtQkdgIiQBzrJN+8UZvkykYDDk45IrkrjTytNnmhiQxEDsnxvLok2FLoPBWVTu7+3Aqn+qY
yurwJbz3hQcLpWUM6abLN3S426iZaBs0oUS+/OdDEMFUywAzKsswPXftmVHEhFcpgpMxRGywc7Mn
+m7o1gIQRXG7s/S4rPvHLAjR6SFFyGCS9/NQgN0OyzgCAM85+YQkIydcU9Yu+x65PgtkRqcR6pvf
+g3Ve7bVNEogyHrGOoRwAxmXMOygdvK6SNlE4EytKNfJlHffF4fiq7X6w9nI96MThQdyD+1s87xi
C+6kthJHBlCy3gm7jJ9+kdEsEESJUkn8Y0Ix102NEfziQNB7mVKTEidUPd/OrrZF3lHdd38hI6Xn
Gro+npn7lPAjZ/VXxPN6Bonfz1NgGk0aG2L+/H787lNDIA0H7I/1FqXwZ3HdIbLaOFiYgU7haUOu
jt/3uEnpYXSD6kMBb4D7NOsKQ1EQMr92hwpIyJcrzwPqnnVz5mfBAiK/5RlgfYJ5Rgqr25UKNO5w
Nzj90IYWfWT5EHXnpNQa4GOn93BfQ5/YyqydwiEnTwUQ/MbwUucXaXOomeQuOAtrihrConuaLrgz
EjXh9eD3XMKDPUbgLDsa2gWvh3I0UOAgFcZMQlZwDvaUCjBBqvi354E44pyoHs4XL2Tc2FNokZwP
r8tGft55M+dFnvGXSRv86IAUyO4rv7bdeHSWTLOtBMBTQL+6RMPrukM6VN4GaPGRJWcpIJEHTkNF
c8akAgGLgBso30+8atM/7FcnWPdWaHt686r4t7qJ4F6OVPrn3inSQbPZNhkgd1oMwVevxJBbuwpz
ur72y3gWcSUAqxmFRwzlqOlZLsaOdzEzI2ZorBmr5VUgezDFSYXOiEWZ8f1p9pVnOHbdlH/7TRFU
BYb61O1GjF5jq7zAcjjxr6TWsxnu1VjKLic57Af6wUZhRWLX57PwMQr/a6MHMUARhIw4eXKvrje6
G2IlZNgH68hKPgPOJpC7eb+Za8Lck+SCSi4gGDyA1PfYTGf8i4VXjdlXnPY1xTPXe1XFauDbl0Dx
OVb4jbsNk5qFPfGcDuTvftSHnpysVOthm1k7SqzWcfYfVTZwmjMwiurYS/Ty7CgX1h3moabfirOo
bitib/Q3J3ABHgO/QHYggui+em5L2E7UzIB7wdr4FnzAZWTN3Pdv2c5o7hlk/gg/VIv1m8Bipg3H
CbD6raj7u+8WbgK3Sd9mOQqRwl1EBkjTdmKhjZZhp4oubT9xuXz7a02ISqLjmW/LLNo3onIqk+2M
ZMKcWdO0Ju2wgAB9nmwbDwizWVWFCFCu4QSUA8CRZSaochY4oddsHDiWTpwhFhaeLez2wmRWxIrW
dIqfHRzOkbip8/Y98OQOQVawEDc4GKLW0+h5NZPNQwEQYGQlp0g5CwBAg6EvACXQX3/gGcmEAqKf
Qf2eI6UHwRo2k58lWtCkLTbhYKiYitP0kpI9ionMzR6X/6iitBiZMb9w7FSkufsdC5HDtFOK5tsF
pB8Iqdf4AQ9NP+AMeJ4dsXMJIzgPKlFzG1FWL0USirWOW601Ai9BR9vnbXk++6wM0QVliVEKWquy
strhgMO+VmVpHBt7iY/Sx50ok2jkrDCxKmsXtu0HzwU5UJOuPSDGubWNsK6vNpcCNEJ9ezt1RoAu
wGZobZO3jgRu/72nkhwgXoekLMyGa6K7CCxt1uV+CB+GwkS5vHRx60RYDi/D+30QkZdL0WT/iaWw
knFMMabv9395LBQF8sam24y2yPJRPu7oiokfKwJ5r9YY+KPb8GUFFXsqdm+wWY+uL+qO9HmK6J4+
vIGjq7wUeH0gpU5X6aTHyQlCFJ1QcQsbocnTRYQ2Dk5q/Qv/KMXq2ik/H2AFo/D+6ciHDhe2azd/
9J694xpaQ3FjZDuWQc/Pmf5ZmHXfOGxEKSVF9BDT+IayqtHasNPMGxRzjqe7qszKsaCh/+1nsM75
t5N4yuQ36lDnPI9le3J7KZjg7sov1WyUaao7tDJKaYbiwkXkGOOYsflLgEV0Mf+mmKXufQC3/sSo
TOgPz64TSG8RzGaLDXGlZA3dKJ6UlTLJATlzCcjH3b/fIdvpIDU/RFP2sEqIwuqom2CyAiDg/PDR
9DSVFWxZurhIgjvhhQ+Ypsgd/OW14GQXADlraSeGs3+Ilm1kXVqZcVU43Qqx63WH0KjGS0jml+s3
pZamONF7bcrxpLg+eU3p9tZvAAQR5bicojr0UuG6NDcIH8n9o7gFaVWalVfi3R5+8MyH+s4+sqHi
ml7XtmXMSa6UZpKiojzEPsqU24Z+FzzFZqYGduXX7AzHD+4C7po8CREIxRy64UbaXT0y9Ad4H4Yr
Ib9qdzpjOYytIDw6wpa4XvgMt0dLoJdMoJkDM5sDxg0vlhsPLTLeVOEAOJS5U3k8lQWMjA9l7gt4
gs5r2awe3qS6Jfiw1UO7kEgISiTgHFTXq9I7VcCFfnONr8uMIePXTUah1vEjxIbxQDvDG9ZOOvD5
gYrR6JogM1DYZa6Zp+ek9EJ8DX3MFBEJ4ZteL7L6ib5cGlv5Jqy2fvKrDcXC3Hs1y60gPzjBBXpM
bKy4mq4TdsTkWyhHn59hI0YUQI15NVfNSfUycNWEYvUQtMxXDsNIJuqzZHXOtWhhTgocfRvMhOd8
UfVtvGLkuS2WaROHribbNSYsqxdDQYtuMRYwR+xvbNQ/2xZncWwS8sVz1I8sboGMQJAdKLS/dF0N
O3s3HfyegY5uv/fOzWNBsh7jZkkG/3BfZqxzBIdTmvKE+LOYfj+2mGR6w32V4l+4PtvZ0slWSs4Z
5iuWciM6FLCNYd4/rJ4kQsJ9bF0H6ruZQNiwr5A/5d6iT3MmUahA3AYIadcv/PVJijzB39JS3O/R
MXuebVgmpcyflX+GJpptJssPpB8U/3HuPw5PDtypnaOds1eJMMB+/DVNq71E6AJLwuopxO/FS7/t
G1Hx1KoSUsILvZiMxLvqJjewCcwMMfReiy8qKkURBlSOwRd0fNuBMepjW3bJo5mJ5wE3PUDiqoms
+Ob/YyA6xM9qE2t6vgsuC6uzeI+YYYDWpXZANQbqSCvpEk1m331+8Z8ZRqvdfsufe6MnM7G4HIEp
yLH5Vtz/KXF7wtE4ljwNgz/UYk5M78fUBRCsLXAZnuNT7jyuDr1Xmj+nWfk/ICbnwjJCW4kqZySF
/ULSnIhd4vX0pHBGHI5m2wGqCDLmHfL1VTDi9imf+AVi6xndhJFblJXwyN1jR4r94sweTORftofm
C+3gnUyIFS3Z62if0Bsve9yiVDVkZ9NtYyqqd/MfNMyPnUfrsGw+pW+E0VK7mV2TceiLDbA2UbD/
lcOk0GQVQUs9g1uFqlIJPLrsHtkpw0K3fn9kQ9gQBm7vBKMCxvkJdwOl9I2VQrFybYLyNb33kglj
1yj7aRlT8OTTrHLO7/CGGhZjFEtEU9c9ctVbiRa99yfW/C+bbA53GxRUnNaV3BcmbvOGX3C2Wq0O
86BdvI1GZR2L458owZPXiUGzAXJGdgLttxCPZrY1MPTIahTfAQ1xuhFZBdHeOg9jpognPU0kviGh
vAVg1XUIInH9ysPHdtMrbrsb3djmznZZTohbxyCkXUflaOa1bGxQI33pSd2Fp9oCKtK7MhMLQD+N
HqmCDhiSwOQric5V6YLL8gasYz9/00QxVlhcQPSZ9eH13wc280pqDC5xmQ8zn9vHMiNNGdHUstnZ
k/odcclRZfaq6rN9yD/lL+oD2J51pPQofjF6DRn9KwATlBbtNJ80JePQwdpQy8lezPP2g42QwtEd
TYM1pzLY9SuL7QYGcE6rFDjQxIO/AsVE/VTaB7rYU717AE7GYkMbDSr1nZLAssSNR/EOQVfl33gs
d54CtN8Mn7086NWGCV36YOzDxdqqS395yByn8L0ZATSRV83dAviaTCQu2T2R4m0UvODuPg3v8Yga
lirZ0qQwEmhe5V4pft1lim1czZcwMnO2AMKKP+3r8GyTe8tZTsOXivcZLiTjl9Uz/VF7kGrBs0yx
5Rp/RWjL40F1qbs65dNBvmn7e1QYMvsrKQDxxfhRFchG+xNxkZALECbHWzm2PFbqI7ybWuMtwK6a
5SgxvqXPYKtwHKHVX8yYmAndzqLegOntvybpAQYNuvVZOR2UseBkZYSXFIj5hLUjRv+IF2nPXHS1
Huygt7Z+5k7bppiHhuu1ulaGZ+V8aMuNtOaNz1sLIpEgckfSf4XsdKWKG8VoazQyWfLBYquMmLxK
ca6AfaTfSyFwJyUCjfLoZs7E2Yu3Wwp4Qlg/7EpsbWpRopQFOwghgrmAXV+ZPSL0YRVKgCrP4XmG
53gKMH15aMWqWt54+KEPCpdcZEjhrTDKW9iYaUKT2ZC6IRQuuk8HvbQ+Oo/mZs+rdOO/nEiJ4uS9
7wkhs6PFKS5wt9svXzpLiFAnbaHJ8h3vIypKsiwGl9sg69fEfn3MdTT6rWXExW6Bt7q6nQuLpk1O
PgsSemptTS2mYNosdXkV7ZBhKDRXC9w3OcdZrNSEVjSpzsfIZhrMJn5nuf0f8nmtbfUdfFXulVsd
cZVNnV/1A+n4FbLMwprzfdtaNK83M8yf6SNCbPjV4/gvZVKO7ACbsx5FGg8EXXbYt554nuuHtfl5
7E0gujsLDWuo1R2N9bJRwMOsoJKn0SGGxOZOwERCfabork2xtD59JGsxd7aCnZFPk5ziQLb79pOV
gH+RemtPn33U6m4qo6qNlCjEND7nH1WVSiOKFlQys2HAZz5F5c1iojEvgme8IGYmMU+4UKkHUYFo
D994HuTo+KMyd7VmpvkMRHVMg7Rk2kdz6pRmyYBizv9hY4i86CVcFnU3+IZ9YNR8ytncJ96l5CqB
g390/AHNYMkSeOoPl7G2PBKeFpAxqyFNKdLhc53j6H/D5N8qCb+o7YbW4+fqbEtwAp0yYytZKnVJ
GiEWHccyw14y7bJWaeqi2uiAGQtrVxeqEtuVUJ75Nbm4KYfOD8CLatTovd7D59pJWxPrixYm5dZW
Xhukxq35DW/re96l85wRHJsv4EWXKVnYxdMSFirmgChm6bTeKTl6Pp5WHrR/haffpbCffZ/mA/7P
mxIE5Rs0aS3IroTipwKL00+pFqXYbWt/5cuW0+dZdiJGPHMpgow3ZaNZsnN3omqMcVown0sL0igW
4h9UP5mpMhvb3/NqD7dWRfYswlDhKLOtCzMjWQ7OX6AVLavXqBR83Lyf2QVX6W3tsoTnxCUpd1td
8IB1NDisK13glfWSyBYu8NRm1Rsk1iUEBFj2G9X9Lrk3k+6ZNNSEzu1baDIJUx1OqpZh87xEtsnf
dxgOJvfmkH0aD1KmieG7LjMJ2aRRApyJlEKuL1MJ0YrK4dfrELkenoq4j0BJwUOZP7wDzX/og6rh
Irjk5BmdtV8lU55F9KwIq72MnE9DsElpHS+gvdy3lxgbgfcqyjvJZ8Mne3PHdU4vdNYS4zdYyCk8
snq6DmLAF085UVUZ6ZeqbAcqCf/Jp4aQxZ0cVTUtXXVdUIKdh582fWBA5I0cqYrjv1ipUqvHMTHv
dp0ZAfhrQ1nidNowg+Ay0QKDJUnCZZUaHibFeUvlV7J4SiLR9Cpnt0FOZmBuYLADfxie0sovwuD/
2A2nAaBYE4B0oelE3HB1Lx89H/Vy6IJUMDhvWtOuu+oGRvoJDTCIrCq+gOkURAy/HyUVASJLhf+b
HEhi1KhvIDDm673dFYMwOFeFma41YES74yBOn7126pRXhEil7wIz87GWN+FWh/jkTR2h8+k17Awd
h4Nxa6VinrJC2FrIImNfK/wIkjrZTxUAj9OVft+jt8jVB7OyusF3kykUOdtHM5F6dmea3SPCoIEf
nUqemqKkelRbhRw2Y8LOiBN1mzObvDjoAyMUNLUL0AJ6cIFDwqNNdujn7q5fTN7OSEI3fh1CYLMp
Rs9S7JvjevhbIBHN1zv+UCUvUWKJR3gfuHIcnAltHz9QqvqQrm/PQekf07SMXcGaEbBjgL8XLMNe
ODRmnPmL5YiPaLAZTZltUIZMxxl56f50kanMC3lY0Jq4pHhz9nwx7KRefEiuLdU/iigtKEm9b5vB
8VjhqzeRcMeU8EG2MkCTyH1a7f1X8WSANcoFHD26ftcv8+N6+OKN3HTFoPsacb64APaV7I7iV3G7
CEn4SF0Bn0bdSUbShGw9mkWYmBq/b0giT8K1Mg5XWThs3v7aagFdTqM9hESpU7Ea9iBeii6dzb/M
uB1k6NtrRa31eANXOwwfqjPZVuo2YVAdE2xHCd3kh4E2BDasSnqsgB4bq1TJO9dkcAfe9G/xS9j4
oT1EfcLe3aEQNWu0iueC1kV79lSZ4dS0qowPWre/RQcHouKhZkStv685ci/ThQr5iaHlynvPNaz6
HF5sKxPFnj6LBQ+1+fNxDgn4iIPA7pk31MPOAFlS3sNsCQXZLzod1u3FpYdhG9UpYNrB7nehHuEO
px65+p2NOi/5i5rftoPSNPRJS2wooVDywodVsIo7w4apOYImqO9WdAMAPmbZWfDaYmlsIwWygSZU
oKHztli7CCcOaM7OLs/rNrx/spKaShBOTJQ/0ChozRQWftRZ18qdMJRm/9ymWnNuxUT8wzoJAv5m
QZwiIhN06m7xA/nlHdxhOyJiWJGxokGpLO9LpsulLKhXPpA+3JzUDtm7+HXeGIW5FF/Rit/0q8cz
qRYXV7YtA/5RQYnVCCgxzYrvmDZb56yBSc50co8JRUiz46psxVt/UTXrFj2JzvAbaVZWbE5bhkLU
aIU+oFd/NCGGU8GDv/9xjdpgBYPSshO+4nS+oR7Pu5GUEwYzQjYzhc/Nl+/zOtTwkhk+0+VhYlas
FCKojsxJKL0RkZqhaiMX0x8raGAo0tBKWtwcjwEjPcL9Cnj4jrODdqLdq08bCf5bJaocYtWksFOO
WxAxBfb2vi7KTithb7lAwez2shGsylvBH73EXzDR/EpyKFW7LbW04vr1WShj/qiDN2Rt/OlOqUcf
gNu7a++tS5P0EGZisUpbz9mLfmCpqNN3XbMRwY6Xk2/FWuF0WwrdQaEMKG1N6SSh0XJgY1Ho0drK
cszx7LjJ8keeeQ1Md/yDaZVddMYBsjSnzBQo6MoYiL5RKXa2j2QgEErn0p4HyiOUZb2M/TGE4OjH
9IdgDQe4BXkq1gA0usKO6wdfeV96ttiVwZXog2eF1lnesguBuSd/f54bx/L5pc7Xvwo2yPIMI8hs
prW+8N5MMQciIOjivzdr05H+JNwX+dxaFG0rbdGYvDxhZa5QGAicd7ZAbgSMILVchJXCDWfqH9ZB
FQZn0KgjIzVru/uW0fk5mlqUdIPAHx9j3cMZ0idUeqgm8HMNCzX7hj1XPaONRa5wW5UMBve8SiBj
ga5detOmNgz6c+fv13DQSpnwov1UzDZCAPWlkAdsCBRpSVgtY5+aA0XxuIWIHMcuL6VM63BeHvS7
t8l5p5CxohCuIEXvzBo4AeOz0Xyl4h0UkQpeUKqQBDI6PiLz9PypGnUEm6PDlN/AGHIXkR5QRQh8
we1jr+b+L9aAScRbcWZEmAm7v0G1i0mEnQTEN/98Yc5mUEg8df6iNAqnazW05bdLKeSLv2lHBwY5
xxpzkWk8LFCQYSomTt1mj0iKE5g1mNFleT2YJt3iMsadPCpUqx1GNRC/DYEH21DK3Uq5wGvY3vKi
YBleFCXjRUNxwRlvlOzwzPLwG0uXQsCufWcT6HDPKN5ijbTwiRVLqGtGzHsW6a6v1EU3h/LltURv
Jvh2/sFoMFaK5p5SogGZnpVE3cUxl4KgISAb6CsBnl+0vf5Eb1b4BUN+ngBXsAOJcRk383NCxgzN
NQXmSeqlrHa028MMxzKNuKMbZIbLtgEUZ09qVMVCqilVG5j6i3mzvJ420eEroB7m0e5TMN95VTtZ
5wmrRcpJ3bvmZ66cy3rlaPiRvpYdERHnUoGb156y4xM4LdXzOKboE7s9lzf6rXoctMZ6+Y073UH+
eI4igJ9jqbiPqyZALyqwJiT8LHF3RVP59BhsBxzxADz3v5bfQsObhPbBxEmIJG/RhEsLENFe3TdP
EAK3SZUW9uu3ZdLIfiyU/Dt/EASXxTTd21GZK4CuRA9WCi+9oqB4kzJFoO/yUUT6Qz44E7VyiJiM
NoVljqDtINoLmyCyLvu/gd/MgxFEJG6IacZwf7B78kCZrf00xboDcYCBEqqzKoAiQqt/wl+3rKE+
JQKA8dbh32qCCrrGctaMVaytQPspYvXoYesd6+U8Rcp99I7eeqS5i6yF3/1J7AWWA5217S0elHze
UpvpvYaG8ZFLg0Md5cdM6SCTSgl8Kcc5vsqt6HUcaUYFPnEUqgOJxRwkr3hyoWwI0u57RF2gm8cA
wX0UkMCzTS1GGwnksjkxOgNKI4fRvNM9VHjHOlcjE6pYy3eOiE361AEy5MteCnDnZwPbzctdNWxg
7itK/yDNP7bSPvWyDZc311nJIHnTzlbEDisns5iy8uu0akKjHldp197tErJd/2UVIAbi/cuaPIgo
hf+pLxfNVDSE00hdWhx2MPnwZbwuhUBD9wuqDwpT5w+33MNYMsWf1XiN0pSVSrAjVKIoYDc1QXeV
l/YHCAzwjLMzO6Z1gw9oTqyr3AyO4keVmJrhTNYETpWUn0oYlLfP8g6v8f8ZL2mJk2hYKe0ju/3X
IdaAHGl9LfbjF9kqq7re+whWdGHtqt8FjznS8t8z/Cd/FglChR5C0omtelUj+rE8c8nW/qMUoi2E
YT3uqpqp9eZdeQYR/U/YRHAyicTx2KU1Y+MWPOrPFNisrsAlbytXtnqxnFZxgPlaI+Bp4tQw9hq9
FdXIsC14CuiNiwSRRLM9hsr8rShl/CDVsK5tNtuFveEnXWvz/VfJyLDtIqGvj4if1bRzGyztO0pn
4N/uj9+Ws7RMSkAk/3qHKfr+AYnnUgoOTwQcPOHrzo5Iq1A/ZaEDmba07Jz5YTHHYBGgeD/eQLtU
+cMBxtRB1zwRvUu7et/UnoUMPAY5NYco46Sw+eyTEBnYLGuIteFGODF4x0cIIe1fs0agGb7/2FRv
/cvfhS27UN8VB/LPKiGqcjs01jBV+peSycDnbpaOCS2STNLFAQOVim5dJaHco6iKwFyNbNcLrgv5
67XKkFB0qz7UPufOrwJP79NYhjGQhovS/QdbSftv8DhSWu4PF492CArOBIdNbcFYeOk2qTmV+Mho
8fvN0JZs0H8dU7f23iyClTRwbUgUrUkWr5ENOvVPPJlUEKKQdvxlowJQ/+CaAqKvbLi4ZB1e1PiM
LzvzFZqyBY0t/FdWcRvKA0ne1MRgmXxo68pYbQF2o30cTofub6W4jM8IYGCIkE/xy5oL044J/eEj
Kh9MyfbL02Ft7z6YxNVjtujEzWJvbcpXmX+QlV+kgVAxc7ArqMaGfVEDcTHg8WlkMzcA+pPuejPE
bPPtn65eR1+BNKg/ZmwtYjYKQPOz/lIepibPInm+j4lD5ZBZAJICgbTm+qsJ+KZ3ydXqNxM66meY
2h6C4o7LKSmO6s3nK8MxPaxavqbPfjSU0pj8EYkVl3FQL6x/6edasW08PZXdhKz8fIMg+6EN4G75
08pG/rHybB+Vhb6PUNYuq6b8BVHimLSaTKOUVRVcE82Dr90N5nChGjoW1C7ECWLBImrn914b19Ha
cUIi1+pniZIiWCCh62G3brEzKB5S0N9vF2QdpZP2jwYfv5FUJW1fH80bCP2apoKSyQjK0gscavpW
+7AGV8s/tAYMYk+nVQmYU/eH3B8ZwkebQn7sIX6IBzfCQ2mYZjeDa+Hz/vdkTIB7Laxy6t/23rsb
fxLBY/ni3dro9PL9eGXp4qSfSvuvXgBmWT7vigJ+8hIAQJ/vhGG2B3zS1rEBgpzheoWm01R4yjSb
J+LBcqFNR1wqlEpLa8RqmgQn2rD6BRBplpBINKn+hX9VOAlnMndbZRpBCJmS8GryaWKJAATtnXHG
n6mclQJX9C6PuaylrH9XQ3RPHiI7nYK2B/eL9qSwXLR7jPN9ZbGyEaMtWhxJDuNF8Oj8cwUVy14E
kxmUFb0Iy80DpgJTbYobKuOfdGKGhSN0Ra89edbCDVRMVmi8IplDCHsLsAJ7iP4j5LDWYgDi4b2P
QECsEZZoNtyUs/OUExXDN8oGLJU8yiK7eHMQd+cEH9qFHRHta5cicoLcFwZRHusctSLJKwx2kuEA
DEY6fi8gPFaYGoCaGL/XgwSTz9/VaDkDyrgdctSRU9sBPddtQOtIlWRjYvOvER9usKzkcOk83hW9
zi7xqIwHwVRdRbc94IIgsj8T0+sKuOfpAhfTUZHRQlRwrydelDS5vkt6Ha/og1H0UphuAugeFbYI
O1fiw2/FQdHBB1cTP/ypAJTDF5/T1U6NjI2Sy65DaedkZWaejZMZBYtaeyvAsw9KxM7mJNt2O8+g
cspB3nXOP80EkPpFQXmMrbsuyKsn+aGp7uQaJndjMhsZVcbR2NgerypzpGVOLOooQLFhV11zGMs8
zgLa9IFZ/sQ7TjWsGdiDZ/a8fo6aMZ67mlY830I5RyVqpWNPYTYOeebNFgzwUxGBk1huWZ3kPVQc
I9l1yhX7/2ARvUxoJlN8B49nRN8lM0+5RTgdYjR91wdDKXnjOkyar/Si/MejVjZbZiaX4ZHvX6r8
OhXflWNb/EkQVZNX57xG66BrcSFkil9h+8YcO0FJJQH3hOGEqjcBFYo2pPxCLkUmawhOj+42+uzS
MB8IB41xp8gDVQmHiE4Qszjat5oPeGoS4E8QwBkfIINUFL0yb/+gmWnPnX2WkDHUBLuXoZkpc/Qa
iVun7iNY+1uKW4r8c5KXWJeqmzZWfjpJuIS5FT2AW8Ib9olAyqd3cb+s176amY7GVlVdYxy5ov8i
SJupWmI62G4NXiqBHK6xWx2ELxZ//bvJ3f4JNrYkEqUiT/RJe0cSn9BM8YRYugU1n8bGdPPA8nCp
vE8PLcXDIEre7wfmvzcIDSyJjk5iw+whC8rL/izynVdiVpOKOK2lURZNzsE373MW6NJcs92K/mWr
tkEFjateM0CNcUqlNPZ7O4/GM4UIJdBhJYIo3al545/7By9DUHZILsJcfH+dWSuzT0jzEXjT/wMZ
kwzGtQZe5J9EQgNSlcFCp9geKvea5fKVXPLpV6+JYfQ92DA4vZNLpxrxzvXxLi71yq9j8lBxODmM
hTckhvgfYUT7MbEm3305kmJD7KlFjqyvZKcXlzfehFjn40qJznM0HdGf6+IPVIOpfaeZEkw05SG/
H0fDv6n4KCbSE5LIHHHRh0e1HJdGHmMaaiLIHkSmcIc0nBeG4PYH5qrGvA8t/wtfhlR5Ujiaaodt
+hPBlnbyG1HFtZcdnVbI/D6OssCvEoHoxJoaXqXez/sxZUo2n2hWURPJ9DqVBkCPbv+uIUomWSXW
g85umpHE1wzPQoMOvqtVGSzaqL3h17vHvmA0T6RaMahhMs8O4JClHHJnrSLpJmi6olCU5+paCiB0
zqNPtA37zcjAJr8Oxmdg651NiWlMfquTTllqSXgQ0K+gtCtE/7xkwjZNCn5UvYZEvC/t9p2a267j
JayLzM0j7hZLsj/ZR50YYhrJPkLt0Im1AUIuG0+kqltbbpPfdImlquU52FY67zaWRn8A8iTpTuU8
/p85LP0eA14+aIki9XVO7eIwl8ccXT/RLucFV01caRuP04sLCAMl6tOBWm0u5iFdpvqV87IUmi9F
HTNsHO5z0A/sbOeDrfY5QqOQEkYgBuDDkP7uqUh1PP+RUJv8fk8eSuhdMKeIDyErW2gbJb+YykTf
mjnQzqp3IlSSqEDCTeZCvVcdwmFO/iMKIlqUpyN+f2TA79xKrMbyaLnwDvjMX6faxBXXvOAcbceX
jTAYD9x5R+jz6OmtIMxmRs2VkFO13MM+cZlM3gSBTHLB1Fnb9PcnlzGKnGVI3Tqp7tBgrNTSGf7F
tfPqm7gXJkwzAn+GISxR0tJYkqs9u35eBHaqMd4Iovj08bYVYZ5yE/GsE3ofCs3Qd26vZpxCRQwl
ODSpOOjJ/472dONqwpfgDmByZjhiS6Jlhy58Yh6wirl1F9+J01xyXYOOGhR9U6eBljZpz43+ae7P
eWOBj4zjUUyoVCKKwfdXO0OcDJEtFK923pWn4baKeVSB2FTNha4nbPI50RCGZUcvYHp3M3e49+0v
N3M7ycUH7FZpTHUDBQ2V3DZ11QGCf7NSMKijQlukPCHe1ECU4gbPSihVFvFVs/WLomkfYwQAuEMo
nR5Sa8zuVTHMImhTNiwJJYzuoRiPRmeS2S46xMMqdct8JC8ZIW5oiVlEiGQb37Hn0vDKz023nuVz
qnyFaHwoqHaZZ/a9WHzut7tsj5ENYWnDGSGSa6gIhlZi+smy3+LJBzLdT/JzCse5iR9OX1VbqulP
9CKqsgBQMSJXoRTtwyzTk3XMzdnQFS0/Jx8g5q6zRtcWowGYbrEKokOx7v1XQsdqx/BaDAuvWT76
603+48oosTegk6U1vXvTYtpOToRBS4DHe+GplZw8eNZetSE+VsV9hO94snTMqqp0LmSmnWAc6GyC
KweWRx6dWHYW3AWBor4C5hGLsDDdhKhEKLGX40KyluPF0+Er7kXeGD+A4lIMfbmvgjFOmva/Q0zJ
DmJh08SXfEXvgGrZudtrFwOQ/vmjWAnt0mBjicwI0aibSRHT1xKRSJOpFS5we2ZBQPADJE4X5mK8
DdnSGSocdNZbFw8fqSfsNW10sNstpxQAKSHwHgbklEc6VZUbmLM/a7H6M5gEZgW9EdS5KwjbzGny
n4y3B943FV1JyI6H2dKkXTWgfnKak4Ck6S3fwF/nnG8+fpwSXfF26Xxqu/Sl9+dYEuhh22xd6e3G
53TNKtDgIbyju9NAWPTkI6mmQA6lvPsPuMvrtZTGDIokKgcODppDVT8C4vYLu91NF6l4cwx70bpC
18EyEWu4TK5jLgVnnDffkXGFyvcv5y0+G+q0pl5LXOCCt2CHEMOVJIKjQTz3YWBpI2ExDBF0vhx6
aq+hZlcZIDEI6H55uj6QBtqfycl7AFji4zzLoUMC/bqz03/Hg1FwD5/M2w50Iu/lHp3e64BDQ2ay
cUv2h73BeBI6Zbdmzou1/aCQ3QDZtx+0fwsh8obmVcs8L3fAz6HOKHeuglDQ/RDus3URshQDTwzf
TID4ODN5NvTqZFGjIB9Bhk7ZU/0leLb6DcvetoOrMuv7Z4zAyc3zKJBiAureyzGQEIchez/Zu9zL
ssJtKr2aH8vN9+l77TZ0ZUWGvOYtoKbY2A6PCPYqIcOrPZD0BkEVeFiHwxVeeE8HiKVcHzMUSCLQ
AJ8aLVcp6bTWNcUxy5u3g748B60xxP/ai8qREc4eW8nOXvHhjRCLcB7Lyn3nBDHI7x+S5g1iOT50
nw5M6/GRgGnqqlr1/7BJXGrmpXK/qL+r+Yd9gJgbQVC+Iz/vZ2m59/y9qCYQDwBVhgIIOFG9duri
70p17yvLwNEs4qjZKytWrvaz1EIczzK8qU9H6+CrSmg3rwzg4zKVyhN1lFKfrwm0CIfsO2GjoYGo
L2w1vWGuAlWI0TyBtOhG/Vsmp4g97OsXiFRnah1kiZPe9IUQ9C/zNkVAwSzxPsvMBFuazEijwe6A
ywhwKeF4yM6BCxIl+DgF3WmdOBXOP2MX9csLDUEowHNX/t2HJt4kZs7+IOwPe4QFKUT0pqe1z1IY
wQN5gD6+WKkNPztB3OLN+fh/vDbvv8QNqzMXItQQxVrHInGWU6Z0YLmPFdkNtXpwErg1t2sNjptk
xgiKkLruN84hA+9P18lyNzhnpjMu53GTXRCv1hgBFqpDfCU6PP6C8MIFh0PrOMeyklZPTj5MhOOn
2y5h8Fpiu6NA5ZxBx9dSIzhDfMg9Lum4fDc2aKKwYWgW58nBoz0ZdW1luBycS6gCdtUANq5ll5WV
zLKVJp56izpHderHXTM1dGpYyxIu1Ppy6U4Xg3D6J+vnp/LHShAo0Yyux8vDWEg9Xrq/dqJKL/9D
DFBK5s9OgyUFXrvCDHrXSyAov+cseiWNwHXUZ6hXFcY6NHUrT+TwNEntxOR6Lldtk1n1ApvzRo9K
VKy9IaX8dgvdPENF7tpVhbUXgwIxR7uvF5pn4NVgSiH/Kt9YH4pwF3MebyT/I1D0Lf4qgbkRed1y
hx+5al1LfiqWRhSMBR643AzkgE7POlYLY1brmKVfuWuUzHwjE+yVLB5SDFen0EdUZ/wsndrHwynO
+YKRf/CDzTuwkvzHYtrYN/mrjlA/tUDDxiijQFFGOyF+E/KPo0aKyqka0wg+Xdh85oAZeHcDjW8j
GpIb5Acc7XZ7cfJu3VR+lR0yUpkAA8WWtwGz+ot+AwsqPgzNSfGNwdGlBniBEtQyNlLlxdS2yxIG
dg0xszSTKFVzAOXHDapWtDc2OvCBREpBkyqvNGd4dPKrxearXDQIlbUYhKuZ/6Bv2su2LQh5ZrwK
xCqeet2z+D/qbtoyAppoyUAF19hhAAnhMR8fqFHXWJ25WxFA7iCrR74xXIrqFnDijB61cwYWF8NA
IexYKAIUudtMsMeJU2ktvCnT7Sq5EVSDClYRsxZ1UJM3+tw4Mow1MwvCMc31n6TNkmEB2mkmM5bv
tGWADpzGgn94w6ZhUK/VmNv0c12Qm5yYqMX4ht+IgaVqoSjbJXY10fVUkuJHGjXcofbUVFNuJT4f
bD1l/NGhRZF9xe0Y01WnSGpt//uK35fmIicdFIAWxfJqpC2NlIOQfU3Dj2OMZqiR7o0eeDXNihn6
1A/rB3sSq++bD6ECwfkHY7BD6NoLaDTkg4Kr+Y6UVUxRv0krK7aPreqHBoAuZ2WrLNCMhTbd89rn
45DNkOW7DMJE5eNivCLt8p0lQFgBqtpY1lGHZqzvEgOaVjf1W2xNLj6zUXSEHZZyftxynGE6i+Yw
tBiNohn465EVOBcgwNikJY6Z02G4MkiTjXC3Xa33IrSkxDvyoMsL4D4U8IBnF928uuP0zpyElvVI
KnBeRgM+DyUk6wqqgVhnSQPSZ/ahB2bjQj0OfJKXgoKPb7xdVSrkLja2/NBDL9w2n1iDoC6WVZag
0JNZXPUwFvf2B7P+Ub4ActCupL0fQJAeLWY9iUfDokfKCMozKaHP8lbkjesW6w2Kbz1w2mUQ7MdM
Kldh+0FEKYQvjLpHmNji2Ajp+rWFG0FTAJTn4ndgR4REmzAFHmIR3dFUGIMn4yaRq35Rf2U3WNAE
NUICH2AsBqYk7Ij0oFaamIyJPNerCOQN0Vv++V+MoNUKIZTfA2luXGA0QuzQYLnFx0bwzpRK71i4
0GUhEZlakhDnJCZ0T5OgGSFxwXrPr9rAAzppwCxBcAcdaS5gpXE0JKl+NmvceFru/hWEIhlC4G/D
3vqw5LS8mYXOUqCddp6YxMIN68tlyqEnj6fZfuLFCwF20fKymAp6q8SA1ceMY3+W3HuARucTB4Ep
IX7ktcT1OkAdiNCA4dzWjrnuWVjxpEFjhxU1kZyuJ4HmwdpFlkvMop6u2MNKuobalU4TTpiPJyDH
n/a/d1taahLxhkAYoV/OnIlZoBmBuIrnwt2W8qEpkQoDphKzIKDskXa8uMNe+jXbwy2OhKuNWTL0
lO1UYyfnlhyEQBKXjk+hhDzhxVK3xiQL20WicWikIgt42wZ/L8DKUMsvsyxDecgt3sn7vMmaN1cN
L9A9oziGaITtMNXzqvB1qtb86SSoq1qaSGZh/nZHSQLsROMM8LUJJLmXtJG4z7ttbxIsKACGBemF
dEtH0ZN40u+9N+JhY0Uk9llaHAWxeVqf7vdDjhniUpZWiCPP1DIglAG1gYbYq/pIsqqVX9uYatgp
LfAkaiS2pa0iOcR2yMYa4xrfeD1+hPmnAGXJ7QZXNH1l0O6RQhZTFrvgiAGA14PrYI1hvygmNmg3
jtxaw6M691zbKu7oOq34CXiAnjU8v5Wor1YhLIcYLFkIW3F5QZfi1SWjBONYbiuCLj/YLnr35qQ4
vAcS7auZf+9d0kv+zeWg2Nl7/9vwqtI90Smczem88UwRN9olTkK/zX8pmosdg9aFBOMrT8mfQqT0
4aBSUxYXOqYRmJcnjuy2D19lYD4dqG4BiB8KIImS3Ld/eHgjbRxaYUkUNhDXFH4os2SsjBXhr1Yv
1VvlZVqzvH9Y1mgUUrtlDcDi91EEDinT6ysYrcKk79pog7dtWkzuyW2FoSPtdO/rOHP0uDWIeNce
qhztbc+K8PcWnFHMF52Q2xHAy24BmSc9TJOVxHo+ZsA87scpHzUaSlxcNgcgdT+e4AO0zYvmvHIv
/l/bX7/+safDztZZ4DQg/GwLiFnVDEV8bYGX0zII4joyCVSRQpgtM3ZHh039pAL3niPp2G3tEkUu
BQXHRByEMwaERS2ie6VSI5MGwmkgVqPxsXYJ3shMQulOsKUEU22mkPBYN8+2RdVH9FiXeZdZC3Ja
1ebG/GRQtWm0uOt5v/JbGIqS1X2FuG8MG8yaSd0stzFU3K0B28WFT/aQ+Mg2xBD8TRmJnZPTXSqy
qTKdKEDJBO3Qah6FIITdecbOYYzwo9DAh7peRTJzDTXV+7HmkQ+Xs0gtJtN6Gx5ByKd+0qJw+unY
KETYIWXoQ1KtC1SeJOjkHwJslE0hzAxxjddXYdt72ORuFrAOXpwVHnKFBC1OeWfsJeJMV7Lpq+8V
vH1JlLERuIR9K9IP8JxlA2+AMAnYeXTSxlBgqD82ycAV9xpLmPsFVa2zlR5Z7NYTSxbIAXYL0rI6
EYyk6/tEtG9JMnb2XwZH5bXSkIXzh9xRfXahUPJbjcjkijhy047UxuoLVuiIJurEC7HRjd/OH1wo
2NaL8MccnkeXq8q5iczOtmwtVm8JSIV5vF/uSmgE9D86KjZh5qckZjg55W+UftUmiM4m7eOLaV/U
6HUiAjB3bQ5Atm/nfKhfNJ20RV/nuN7YAn34XavRdY5HrSZ6uovKaEHgBAvHOKNdU8ljmcQMdM1J
aKJ4nDV+GjOTJAIlgoGgd/kNY0yBh7Q6nIgEeQbqHg9kNtkN+SPzVUtSaJswtcysuHz7Hgnn0dyU
CRy0I+LBHRCxQXbHQdZz7yNQTs8Dxv+f8SfVFXWTEFSOIDFlDliTR4GjpCLHzaBu9cyWONtmu50H
hCs+rl0fkRt14CwtZahedBC4+iBFILcrIfCEebhl0G9dsRIBKcw9yl8frWtimXkRFtWaQPm0Z13r
mDPrhfq2diElxvND78xH0fsV4itA/Bhngw2LwEJWK4UyTy8NelQ2OCMZxmycidb+8DaTMrFe9Nl6
bWZEbuFnswlIEjXg3xvW214WGcoAZtbP9i/CLWfH8PnQCcpgCBYZq2xi67I3Jfko9faPn5tFNhTH
VYoa03U73FhGL6xSRGi2Dbb5Uk0UxddYCkRy/Vp8yRHnGh3Sw4Sosx3W6xLKmg/NY79pzM82/6vh
hVi70mIETCi0DorwORlcQ9a0rPgyCbieQUTb/7CIjEbnuCgAqiEVwx71FAnxifd9nlRnXa2aorKi
a8wr6WV7jrHCwYt3qaEHEMlQv5+ODRlDpZ7YbeTo60MGKGjhtYee2G0Gqae3i2xrST+jeBl39p/I
XP+aLA2xLSTdc8Am3vqlCHc18WzfzfA8B8RNHnNuGOebn/R774RDmYZ143Bl+l0P2B9rgxgeQZTq
8ehtGi9eMHGBhW3iSf5YqknYjj/DMRyAUJ+QhxRn0B/cWI+z7YUiJFhYZtxFppVSEIP2Y6/sJnGB
UfG4/G0qK0WlzEznMekg+z5LR3D5+LMitByke5cKIX4RD2sJYdwgQlQNAoGj7DGItPHPliiatMUV
vLbdGh1MVp/Uf7N0/f65V3V5qnXl75KU2BKccij1r+OrBFICmwZM4ZOzL96mcLcl77ELrl4LDUWs
vxy3D2YKNXqutxvSU+SQorlj6MgQu2dP+DJACFXqZDTd6sLiftDzvVQLFVhgLxbtLUKP9Mwyg2xM
LlQNlgLINQdir5ISU2mJqs5U59umXkMYqbvz7fA1OOV2fOyr2yJpbwuKtZnjyy9q/Q88k5fHiQ+o
l31bsNNhHNVaZWw8Bb7A4If65VRA+YCRW1T2hmFdFQvco8eO5Gp/skwha8dE3lAzMweniuyIMDYW
rHHmj/Vn7U7Tppg2thknW6tndV2qY3I9PyynIMmpuPnZxWpa8vXhLrEB4/UFIRLUH7QPBnufOIzF
przshHNAaiRQk+oMQ2VY8KDt+KbMP/4gv66YGdllnu8NswZrolSVqLw70tCehgL0m+f/fGv+iRxn
80Ze6uie7D3X+rDTNpQVbog9tXzGAISjbEaNww/BwyIrbCXwnnUgYOLLk88EK6q6JjKNM2Kjg3iR
Q7cXmIo5lkbauqkY53z2cXspdyeOP3x8BwfACY6/r2VQT3MC2sswIiE6DlW6yUzkDae9UcpuYCRy
JgVLoubUZoQfdgEd4OFEOan5x4jKOzfWVb1nVuIXBk59lMBA+8hSJWbV/jNY55JURRdlVsLfwAz0
7NnrwdiYLSwmvQyq6H2hRo4/btWgfGjLjZCbT8HGvad+2HDdtEZpQP+F4aNaVyirzmTokszXh+op
RrLqsge1YumOI/xeuC3PIKQoiyNxbZftyFm5eQJakQcy+xHmFJ1COvEyjWtfkj4U8y3BPpMUdiZf
mCs1tSxoHWfp6uxyS9bCm8qFhs+gEChYwOQnzycRh1u+hys2+ACOx5yuGr81dggXczjkt4MLSYYX
siMNFt8Kb6p9r6rKSOHw8O/frN0PAnByaK1tURrb28Z2tj1jQ+QUZZgqDj3vlLbs/weYjcEUZF1Q
4Pr58wB94GKYwDHSxxdx6KmivPdlli9UG4fSb4lL7Pzkm0p6ahSs/IzBWfE9TpJ6k+DQaKD1q1o+
es/6lim3Te+MPZeobdlsVzKiQS3zTfEhMmxhZzdazVhDLcYSUNDltOwmQFa8+AH1B8fBxa8SkOwm
yfLX7doo/1IoubU3sle1CyGamBqjn8MFmJg5yZC22/ewI9gQ7/e8zOOp4jeHabc4C/MC9KdDaMnh
bc3fZRbdyJUN3LwMotHhCR5AElLDWKHOvCf99Ue9PAAAc/P1tScor/v1cAFRvkCldl5WScEU8GBa
fcDvJ2Y6s7nmdRFC7QbayJ6FmBdbM/1lNGd31m/EqaQQcKkLBallVtmXyddkvRxf2aGQwfypqVPp
EEENAksFXGmQts+atIeQC8ogTq1SFsoLVNuYMY+T7MkoFdwbJKCgaIwdNExzNi69chf5gSegdADz
bNqoRShY8dhjITM75fUnqgffU11ekPxYRFlG6aidPWHJ04ugZcTHrBdt3T5b2/rKN8ocAnn/Y/0Q
lefFjndcck43bNSJWTR21/y9yEvzqlBHpLOyssz46WlpTzM5F8IORtpbMm0+aEYWJiuwxeMKfBwU
g1Wn7RJlP9xi7FMUrJeG4/1JgWuGa25s7YcRyl3Tr1bKgVZeSOWzSrcbaNLrkPwiYNOt6zbDiL5x
Rx2CYLqtiliaGngHOOrW+NQMJH+PbG5udhUt1/X6DdVmNC65pZli1r3jsGlf/jLJjG4pTyBQyJJq
+W6UxqUMG0iCraow5VRBTjn3aDwC5Kg5O4uPcPonVpEVuc1rNUjBdofhffNQsrixj13Ghjdi5uFh
jQPAEeDrHQ6Xl3h7Byru/gH6U9OJL/dTdUEyvORi9liU/rM3L4m4CBYGzf3BijAs0pUlSJP84YJv
9+EtC5XMs59axnFgH+V9d9D/9HkT4y9xP2zUJ5J/ZsZJA6QLOzfE9kIvoA3iBW70aQiHxAIUc0zf
8f+keDxkJdipfn/rBD3yL4cgBMcjh/34Gc8kM/sx+pFe5IKJjI3PpnJF00JZZbytncsjcRO+qbh5
XZ5sP2pcJGrRfZ+o1kJkRWbEZMLgcCP3NyhuQEsIj7wq9t/EReIkYtBJjkw34S0OwMUw+C83/QqN
5LRWa/sseaejGGCeZFD0Iasuy60FsIepatroC3ESQFhJxG+joJjCkbeUeiKgjFcYVWz2tyqq1BzF
aXBxrX8JdBqZQxWnlypl6l+KbxVG8IbSp+IM03ICsGXidGWUDw+SNebLintpjAb9Bv2x60IDXriU
BD1wT3xATGU4SfU8GOE2J4KwUyvWQlX+PehjfmJ8KoXkVfNe8Aj4sFQHlpablx3dEmh73qeBLOZm
4X4wycw8V4VCmQNtnSR9FDXCTFb43tqMECV4ELKH5PZq+5Wv8oOFHOGdmnb5442kDZt5xU5cVK6D
ibt+fHJl1kCzwltc5EvC+Yd6UVdvfMqHcqXLRVquYZ9jKUbhFUwCLoPG7+NnJv/JHcwYl8u4ZixD
ZeXmp0RJ5z/TJ5yAdH9dwrwlS22F90YWye+qCHXkpPo9+T+sE7Njx6zuHrwXVp4GKvGPORW+w+ab
c4EHitR4OlScsi0euR0sjn7S3haf+VQ9bkIME7LlZzf6n0HVpEjK1hBnxEI69z6tTd12SMyyyNw4
qzBml6dibn+MSBk8M49mk/sj1ZL00yr0SmsdkbBmYRwVZwMWKiD4nBRsFwMhxjRFSP8ICAX1p4tj
YoIEnMaeqzaSnJBGXlMy35J8fxnE73ACVYytl0usnwSSfZnLqAEpUVb936lzYATXlurtfmV75YIk
tDMQKGnoL7Is6ozSQGcSpDpixkjRayQx8E5T1sbg8hb7F8dFEFsHrz0Vre9RDCYa62bTVOYHycew
Ht4OUlEZ43WKxO9F/nj9OgiGT3jzPufZI1JsCQO1iK23arCRkneN0zDy7tqxSvd/G4LoAUaSng4J
zxBBOjORoFsOsfiOQ0BI/JagnjsvXDvfdijszK3kO2T87tXizCWnhPkQednAG8497KTgRgh9BN7b
s6KSB6c/54F1EvfHuZKPitq0ciEngp02Y/vid359MaqOnZm3bhOqpwtGzGjEYOwfL6J89RWX05aE
+JkN9g6cDXvW2NySu9nmu5we9bwFC3xL8cbXmK6/jkiMyWfP16W+q7vA4rjdfQnzRNBuBKJQ+yKm
0Bn/Fk8a65uwYphohjTzDT08MWhw+E/jPMAwhZzKp/bH/pM47rNBRb+Fy9axD9OVy1sTtLS3uNVe
tgT6k1Wlzc501J41CdVDot/pC8wo6etJRTrdvwhqDm/Hmmx/pd3FJ9SphkBKudOHmbmsv20ezD89
/LzSLJtfgBKB6jK8ZpanYZ1UPS6zZyrI8T2cb/ZJ30cjlQ0yJWA9tFUK7lYz8bIuXzo40RipF3jv
LVi+RkU4BDwQQF7bAANJsZITQSvuLwn9YQxV/Zy/pTsG3lEiMaoJMlaOXI/HWkPOLu8LgsFVCpks
yua5A5xHsENFW6W9u5LZTdncJeG85srj6fwNyVjU8Ehf+kQXCEB8bdSGXNCUmfbMKdGZfK9xUOnp
5rFSnD+UruSKk9HMaP1Q9YnxNE0Td+efZrszX/bFknEtZyWQ2urxx9Hial3XCVE095pUqwpyE4t3
N8FghvBSlkJHDonx80kmrT5zKqFxVHUXU+gVaEBsxlR53Jiem3i/DagN9D6+/1wJ6giJ2bzLj+de
yZQubn8ObSLdIVXJEQQrUQ+Alzir2uqvGYEOpSoJ+LFieYkAiNk7Jr8cv34zgjqQn6KzaOOj2JZv
5xqspy+0ApkNIZWtGYpI0C6p7vMwsjIx0ON1i0NklFAXouNrANPE0sddXC35lcTec7NPEjHC+3EC
hThSP0NUAud7mYKr9JjN8lTpo5WdAO/wTyHwyr0YVVKFY7pYj9yTj0TUvCR51mWkRMAFp5A9nwm6
4AP+DaN6zohYu4OtYVsfuTIFC8emec9vtBm+w5O1yvWRKKhPvLYG040zv9jltiBjGKctflprxqaP
IGaDPz+kg2oIhlEhkFiX4TV9TorV/QZ95t1pZp8J3B+s5sTYJ7GfAZo4Rg6kXNMDhQ321r7kGPgK
cOV9Ax00rk7mOvIR6EYTTnrYwQZhATG3xlv8hHuxa9QcG42THI8NIJ2TwqnO+8rvzOSTOw26kn4c
nP/dslSNU+s7uoAZurT9LisaezaZOm1kshPan+IZfdn434djNETTryHYkWwNcYaFeAlQ50VMhnhE
me3PqDHxJSIxxiA0B9unWJ1Sa+F64+EavyoHMJZp98GG1aOA9kW5UD2spTX4fpZU+T34fqjEqXPu
5/a1QZiDY0aiQoZcHmasu68I0uoO+TaZ7wcbPObJaY5O0svmeOFjoUzLjVNJWalm4o6WNUScY6/4
MhREGxAZt+cToMS70Omszmwa47RNpKd18XeZmy/JD/CjtMY2BpZOoMr+Gi7HSt6O7+IOgK7VnJBy
Y/tM/mqsmSsIZfeYo9JjkwwAFtq96T+TDDlrhEcBlyXkk1n8WyxZ9wqmbY6t16+P4nKp7H0hA11K
FXtKekOqeJDczaRzqaxysG443iV4h5A+ci72BHdE5sFLrrBA6pQHdIBv6kQakjMz3Yz+ieGxQl6P
9s5pkk+UD4Uniu24oB8YzL/Wmq+LaNYliK5ukdiuQk/CY6OesdbLgzNg3ow+mVteSmSqZEX8s/sA
mb3kRxUDwWubZuGnyRAVk69YlTNY0l7pa1EXiHQHXCIXvdB10cZ7u+9TjBUKTic00Rq+Ks+SGhIl
HfyMKByPbuaEYusE0xmVc/HZNJrd4HW4SDJRaAAu+Qr8xdjU5eaZEYym3g/uXm09EEFawHI3LFzF
tFz6jAj16HrzvGX3BOOVHROSo2oyeWj0knJlUEJxsS/J3UTZ6ZpmIp6OBOFETrMa6q3qLC7nC/Ys
kdCwaSoafV8glV5yd8tnZdXlREJuuV/A+D7ngv5e8nueEDMvmp6ujBN9DnxD96F9pxD0jypc6Drf
dga5zaLoIrVz2NFoAwDENgA7lBifp2F1yfFJQbpYOlSHPCoiVk4Zb2f924LqQEoYfR+v421W6K8e
zeEMWam3AQcqEsTfLUHwX5/x6bcVLwHt+z3FB/U5a8Kzopedi/uoG8aZyZVmg4BJKFOZr8UlcfBR
2RDywWxU/w5NDNwsTDadRj8ZxX4s3TsKa4qeg4WDe9vh+/wjoCE4tTr7gnt6y4oglK+IH3DngTYe
5LV2+BxqBbCaz7CNL7BcoA0crNzagIY8gV9KGxjcuiGjlBow8h714j6gAzw8fD/G1zh8Q8PYAq4M
N1P9n72NA1Yg8zbjd91lcxkwGq/VX/39CN2qLwlzFYMK+yKZ6A6cN+48TsK0l0R84PbKTZA1feC/
qnZmN8l4KBSZNYFaY5GjSS0twj4lVBw1V+ofKLhqXY5Y+oWY2Lt0WUdj/hhfPsPqqj5+3iPL2N8C
ptYLENvgTiU3BX9MBlII4HiWp4zfSPuzGN2DstaqgjUCDkIIgdl7+gCPHgltoZxGj9jpcqaqKr1N
dbNNPU4QaDWSoZVWfS4wplH46D3TZ5kSWOgsVuCngH/2bkweAr8vIOX2B4UhF0pcr1haSiSlGbwa
wtWUQe1hICRLihkV1kvHMunVTP6xhSJ44ojmyJK5WdA3Ew2Q9bMTgzR165+AV8OD2ELctIDYfPLA
PVvFGfmzoHfaSyCj8uuEbQGvKm1p8RfIunZ1jQhTD3vgqDbytPRHQfoyUh1NyD9EusFtCYpN0Efj
pm+ptVj2F2TlMktIgVTVreiR4QVK54QO/x8/kszPp1lVL8273h1PY8+ljJPvDC2NwtJxiBNcCFAx
s4TPkzbWQ0soJkrG3aUNalMDWGsMYakAkdWfxaJynhZXn3xYYuGyFZLspbofjIcPhKzXeozHG5l1
JOhlwaChHhYmThFxXOTDQS1b6m4lhfLbLIJxGxvnZzGtEgBiRXwEV8HV+pzaAFsDh41HttrrHBSn
X1adBiwe5wa/C6vtFnHLo6XQpPh2ipufgB/yWI4GC+5LeqCg8RcErzNTECiagSesvuGJV+Ornl7O
8+7KJPkR1q3RaOJIyg4WQbktd0oymplyX3KCd243Bpfv+F6hq+zclE4eVUvW45axnGEtIjQIP0DZ
G8Cw8VHQaab7egVMefIY77MPrA1KACAtGodGIMftJardFYxEsZrDr9tzwf9XZpBlmsm4XAE+fSf6
GauRdzJxTXlrycUx6aW8+yXEV8CnpF6R09O8vDcwPTjQPP9j9/OUe1GVUsmQwSrxMH1WKF/678IZ
89JsesR1BD/zFLaisYf3GkqVvELxH3NPDRZ4AHWcgDGf6sANJ1t+CuvCNqHCt5xzFJxSORfApa5X
0QVgnw7womrLR3uyimRCVbOnLWuF1iIS814257PpJ9tdUYGumRUScHjFsNkTbyPiQ5UCtjhvTopf
n4UMWJiwboWfgmZdrqqctsnCKIManH1WKBWcw2oJdgQkv/ESxg1PVjdyqRksuBXBBgMSngWn+tue
1E4qnS60pUmSB8S/a5wAa4YkFZdiVdkxeFqPTsVwROZLD+gY6no7o4YOdz7pe5Kz9Agb5omvKZT4
5W1YAGScZJB49fz6EGCiiVg3jMzWgvG++H04qI8JyzQ9liWcedMeqlXGIziMbr/fWevNlg7EK075
f/QpQ+uVsvczJsMmzNAjPeMf1/R218UgiPIEfj9b2JTKlgc1yLwFIKERw8eIBpSLAHo+eEr0AEEk
GP/AUPCMRwtOimqEbIUKZRxmM2IR3x6ONzAQj3ufpwNYkBYlaG+nutIb2q9+8cdhjAg4srbOstJN
GUDOan0rwFQMzlDRPFNVE53O41thzqdWPpram/1BT3FWPmKjoX9DlnYj+4Sculaw1iYoTe45eg7h
uQDfdeJ++vWTORmm1dgVAXPHiah/B1gULpDQJZ5hWnDQpnoMoXYz1JcsjRxZ5QggWIsqzPnzClPo
huyM1zYClqFJrIqc5NcmMq0MWqDXxQuKXWqgCMvnXyAhJoTN3v/vMJc1PgH7M961VPZKRT6b8WV+
U5+AO8o4otvKOvxR5Wdk0fwFdqU16Kl2L/oDQNT0/7SzXCWkXi9EST97yw4rgRTZj4YD1oKf4huy
vVWEWGF15/1iXMGa5Y6yiNhtjoTrP7I0FMkO5/HSc69n1170WxHnrLU6KJ+/vA51yzLivKVqKpL/
HbiQDJZ9/+NPWhalVmayFtX/TlOA7t/ZTOMUvqg8SVBUeIaAHhfh8Cv4d/Gh844/ko0DX5ToFQZi
vo8YMxo7e3KRugurafFtTNG88f4j5PuoQsOYBGDGeZoWALEe3zE/StzDEnvmoub7/70UW89L5SrB
Wz60G9ZVgkOl5gINwmBXga/MBwF4AqeSuLZgYnuI9OEXZUx048B2pG1b+7B2RsSilrQe/Pab0hDU
FvtbJMFa0mgoirnenvQMGJfjuFqxCi4H9TVW5eg1FAnml4hrLSt0jNXZkKjWJpOkNl9uTEY3y3EO
vyZd/7jCNJsIaYlxdPyzkomHXgVVwBkVkKixK177zS69JWXBJijAwIH05MIHILmqwHhkYvBD/uBm
67EPbkJ2tAt0WvP5XHveH31QeBBKssbllR126XkUwt1cxsmaYr3CoG9+0YF295BX2Hphaq+cCEEn
mJlAlUNwATqLQIoxKyMMbZYK+VkTdEKQc3OKux6VQbSH1shJ+VTGyRroN+iV5obJFBmVvDohlnH3
tBe6NhSre9wrzJk/oZVh7UV8bTGGpgkn2biJEBIAQi//GXbBYsI8yRkuHZ9bjveSlbIGhb02WVcW
Sumdk9jn23RB5mptX/puBCVvsqc8YWj07RgHkkzZiTCgDouf2mgvi0s8Pe36y7z+K6UgeIDyamK7
bXaOMmEgz5EotjLHuEDOkJe5gKcTNUL5pxiXZ+Nmgef698ADqpptuuRuV6pW2IR94X8HBmh70VOq
dRFuv5w+Luk1mG1Ni+5aBHpwW97Wun1yavuDDnOoXWEGv0pqvVp2ONiaZqd3d3AvA91hLF6zdPxa
SRXa95DXw0Ejrq4D/TEqak8NIYeXaHJlHpHXonGPnViMnHdWikDagkW/3FUpKM8oeirfur25iujo
7RxnzT52OU3s+SORPN4HlvX/q3IGNwOU/wGFD0Cax6t1YVYBwYwnf7ldE87yU77kDfT5Z8509Olr
tU9cDTb6iH5ms7RsIAaM3Mhv1ub8KD6LMifi0BBymaX8hvDysVdAJyBx9eCFr5IoT5byKo8WOKGb
7SDJBAmabXkLonbcx6BXgF+h3JDKSOlpb7TFMGEvmH7NmofoEy9ZxI2AFwBad/8Q2hfvywmPoi/a
rJNaXwUInWgAuk5C4WEIS6qfmDrLFwGrhVYyPmkbR4t9+ozutI0sq6q7HGrcfCVklYZwbB4G36U4
sivPeeVarr02h88M7ZmmCQmjohLx+Gs1mMB8Regf+eSXvlJmX4ShJMZGHcyqCuLQyoxAwn7ZLKCx
bhBvgYu/HfUkGIE1Yy175Q9CIbkbvSc0eDguXw02+35Mw3IobCBuLTMzjxo9n8ohXKIguHvdChZ2
HxGXGX0umMqOauoSrV3urkzsibegY1fh1fPAUFWruSx+aRQ427fGSl2tyHDo9rNuaDxp5Xv1i2ix
2KaZHe/l57PaP8w3gilJwyK5ZaYMqaG1ZocxyoJC+Yv5t35Zb55yBI+9vWYanf/q2LI9ZCfCHUyk
FrLIWgkQdqGKc6++McxUOZ/uZ0Kv2G0U/VAuhj4t6dHXh1nKxsqFDEhPNcs4hl/Oh2K4K531Jjda
mus9Cg0ZI+x87rSI+1fbPDp9tyieAApaN7XTzU0KfRAhWHKJ+nkt0Fj+vWR+c2ymn1KjZoQiK2od
FflA2JkPCOqukev2o/QrsAgZi95BE8LIAx8w6Dqw4cahtlLgXeV/4422PytMP3Fg3UYKCMNlt3oj
X3qqrWkbGXeAj2xcxx3IFAS86ep2S/RsRrtmmRSAAEnyz3UhiYjIPW1p+4iCH4DJ9eSDJDrMagGn
5+9GbkeBoUeyXXSzy0+jMofpIuU/r2b1FpNy7qDGpRR04JHpR/UPYH3+wPhPLhdKoMid0HTOqXIm
jIr1yDfJM4SSokuGkhZSM9vi2HKNjjxgT5FS+rExSQB985No347V4qqhgnpUZ0fcS1BulfxEeFy4
e3W7YzFuYkSRf/dCNBU0hIFKJamJlFvzWUkcfWh3CFI8dAkamg83VN3xHBfMhddxy98GcWNr5Rsx
QPbCduiCxU10D1fCoGotoO/Sc7XPdvVHM7P1o2xqxGkWjZB7vydPIcg8tA+cnKAtRbZl7PtKi3T4
d28qG8EsG1oilZv0zsXGv8s6C0yMQ3tWo7WNoMGl2cXz1DJlmaqZ8VdOPLMcQR9wleGj0mXSLaMb
enKhwSztEjeFvISfTLKSeA9C/1LUZBg0p8OHsdcTH+aHBfs1cw+AOWu9MkF8ewbnxVrXAG3gpL5R
EZAaj1lDJFFnqrtKz6Pruih81xF+e5NNx9ii+uN740C6ZfbBomnUR6+dJO8jEzV4j7Qt+M07yWDH
6EL2yWq0RnQiEMRHR5YR4gv2asZC2VW8ckye8q4+hS0nDqz3FjeYaCbkhe9ruIl/kXl8HK/o53hJ
cMwEfV2kCjeVDR0HPiiuwq1zunf2uorOlQo/USQEf8AKqoIYSW6W4j14p+zf6GBDEd29BZbI8pHX
Xu/sJzlZdsnttVlxeWn4M4yw559iLGSJyFqcT3F+gwQHNVvelwzjEwR19gRHm6tgwwc0lqw4/qwd
THJ/2qo+WSmKD7ik52UNv7nBKEUK+DccQJ27wNcN/4wKZ+iTEtFpbFoT/MtWuxvQrTsXK8smHjsT
RsS+/abOHiaSTa9zai0rtKfK76ot5D5/OC+GP5OUi0UsCC9NDaGKDP0WHY+TWx4VYkbyxH8p7R+R
IbgckOEWF0GQ3AJY1/iPQAOwTBHaTDanSz4F2VrZgmMBqnpid4EsMjJq5qweN9Fn0d/OLKUEOhfp
8TOIeJlwlWjCn48JFv7VhyrL7rdExVOQQEP/tm8L/5EgW/kcnZNQX8RC2rn7+a7DmwjCTsE5IfBt
3UCMhPXQezYR99lwZnUyiEyaB6/Ukq7uNHzbVI/BWPmRReb70bSmUA/0Uba9k89Kkex8cAY6+j2C
b46RTVZRDc3t/KV32faD/L9bU/DwUNrFG5WazWjBG/zH6a5XTQtfEX8ghiJQmxzlpetBrWS673r8
k2qj4jlU0puGJwHyWSoYuBeQD5ETy2Ndo/tK+s8PJXaNjHIHtCsGYQqPRhFmT9f8sw5Ko5TUOm1g
PeJsO9OPNjkCdsUgI02b5xdP/s7lPWqAoymRZ+OaW3xMls8qmJieer09DKM64ZHY02DQRC8sAOjY
bZ2uF3G4WKyQ8MbEg4ZIwZ12hWmIVw4rOCYDqFTu7K6Qdv4nPaE7aFe/tyISJvLt5Yg79pgT7dDQ
NkdynTnzz/Lcl8FSB49KKKSgpQMSigYdgaT0CiSA+ITL3ub2/z2p2OQ+X8XSkjrNf3WbFZhRxHyn
a5XpVWVCIefYdRzfHeGt0m6Fy7JZGJB+usA5jt/fUPaNFTAtpqmDrNsHd8yQha8yiYpCkjExaqDL
z2XdQEUsxfC15+j9geTXK8Ms/alLYRJrIdOu0BlDHv+98qi/wlyEkELWrXzeAYJzTxgxLkJki+p8
CwrHlbiE+Yba8wXJwYWTM5MIdZ/ylbj88kghc6EJy0btXz1/TbwxzKqfwM9wVDKWY9NnBuU9hB2p
sy9yGrgncKA3ZO9LZjRFqljAxdeJnwhpeVHcffTh1CZ752xVJrfMSQX2l0phNKffR2R1f8mYt0cc
KfCW9YROoSYYI+5ZZsRhOdCegWwnUV/adsgPI/TxFOIBDyjlBnXw2gdAkhme6lnOkTF3L1blK55U
BDqLxymnHKb4c8xZT4+N5qAGKMIjfAK8KLEM/rRNbsigTlOFhjd6vTIiSGH3eK/6FY3vysu0ubbw
gcWaYHkXKdBvUEHRZZ7isF63M6Ptf9MdcASZNdhpv5mY7rDLiJAtU5g+sbsOHQJ89dPWjviVTE9Z
NZf0oS1dxic2qO0TSPTHAzXFZaqsmyBx8UNvE+mwk02Zqv+ekT7xg7MoZfFZ9YI9OLmfa9m/2eLZ
m0BAxnmLUogDDFV9hKUqLunGlTWpmSCtKi/xNdpCQPSdxh6I+mEaSII0C4qmBBYIdNnBsPGoDQlK
fa4NtWS+jVbEbzg2LBXrgtEHq/NOOwCPXluDGFBxFruB1kKD6ng1iPCzzqWUX7PQIsEsV1pWIFPi
srjWeukX094azPDZm/IaMsnUYidUNVN5tKGcc2dT3pYNlOY7CcTuShHUKzicr/8Xw/HRp9nFb4q5
aBVnODDXGvFDNFioKxCxsOuHE3SHarpN10ixiNJUxKoPdZklFsHDZ9ZJigHKE8NwYYZ8lMO1bdS9
1WmV2z0RE4wMYt0p1hCQwSWMcuw+im0sKG9zJAZ1lKPUCFdIYihU+iq5or+wORpFqdGVRNkwoLon
GUYJ+mO2gvnY09aIfIjH5ocNfhmvP7emuYUz9AspJc4fi/zvks5iOlMIbokwXjTFwSV3mmskkWB+
n4QFMTH7ctl8yibuGSkCiPUCxBdJGvKFIB1Y374u9dWzlP+LXI2/Nsq5nVnuLtinvRHv5ClDe+ab
zHEEiNrt7BuCzhaNaXW30NuMWkfxVmcx7VTG8dAtHM3/A4kEhuUsjoaaqBk3WQIY6R52pf4OO96o
htJ0crvz0pm9VWIkZTzceQ8zCrq7+v9Cd0EhSwfey4j8heuKja+JhefalafePo4LOBKwPJThtIFm
0TfNSOt4F9IkM6312MSFDBYbEcWGoZtDrzFrI/nx3Yx8IXxDDzGoNMmRBFQxG+F+jskZbaVPms/j
gFziX/drj3p5Amx6mAm2hNgWqQxnZ3p8g7ugKDZIiCVphqW3fV3MP28ZWkLc/R8Qxrpq6lgUqLp4
47v1cdHAxZIqnZI827UHYDlaIxEYGFjbSehHJIeIOPhdgixcJLttp4dCCcDX7L405CPk6ptObRtZ
+xxBWcW9Y1tkFU/CSd8Crr+E/MR6Wj35Ga6BDHKC5X+RY9rzUV8LSZkV3vB+IU2GK1gkviUQ/ery
uwmruWk+MvyU7Lih/3cP1FVCUoIijmXb+wwDy58fstOXgdThYh4UhvFZcjq5hMzILPfuaTq6ZLZM
Op8jusqFIF8LMUgV36QcLWs0EaovQIKBZrzu+uRtOypN+CziVWvCUD8dvj1MAFw4gn6BWDOQxKoX
uSfak21e3OD47xsK5mIO1x0mNXdqXAMXXLefMqa5vLPM2KSl0ljyC5wpGbr+wK6ybWQBQBJrlI1S
0D0vn5Hruj8Sr4yrwWQTffETyNQF+EFRHjhNrCuGZnsmJlv3v+o/Jq06lD1epnE1N7GK0bFjywod
6xnx0tBylVdPKKmZRTs6hZmsEcdjE1j0aN1Qxrsq36JC/Lv581T3GA8xMtdtEu5pH0aFxRBQ7o4s
clq1+/wc131jiL9veesG5rpqSyIzQZLAuAyZrQpHJdhcfCJfyUytnCIs8ae/nOx507/Hr6XJM7fW
YFz95mkvOwStGm5juvZRyCwT1G4+BnwPgnSZvNDt91wc+imsPe44P1l9A9YPcEM1o88EzySJRBd3
U4dZYtqs5ba5LLazsdbPmhOSazvpKzEpoX2HgMmy/+bNMSqM2C/UjM34ujNdvJDfM0RXka5ad9ns
Fsgqy1HM5HW2V2u7+3zXj0DaXZq72NeQwiYvQG1q/Tt0rIYrDP+1srJSWJOptDKtv/4DNh9emNtw
EtZlZM33J6lgtw0JAYZQvovSout9EWFeYwaicai/YBTu4yMqyNR85Yz1Z68zGa9X7Fym3e09ptWG
rdvOEqXI5SZWG/06HlmwEtvJljPvis2i+qUq6xigLCh5+b3Btde4f0EIWcSSd+TDQj4zULK37mKK
1X9gDxH5xw00TlQxozaH18tQMRPqOc/h+z1hjrg7kCXgA6oKZ+LJK0x+WJV8voIB68/5jKbMTEAG
Q4KCC5AX2jxcv3myi1iIdiyYzgjTFPs8Mfu9/T+vh0iGTOM9ChIGO9KBa4Ix30HwFJEBpgKc66XR
1eJ9Koy9I1NY2XNxN//i1UVqjn9CdIc9NhjU9JiCafZ8EbrgVz2opYAm5G7Jd/mN2QaG+S6mRfb+
CagjaDlfkwGc3zlqaAZ6Dy3N/v8SztODxD8D9ijh9SF0veD3FgEpGmUbV129igclz+onV1Qvg137
1npSFqhERS/ofiQobkd7u+yoJTl8A1P/IKZ7q2bJEUofZfZBPvgDVUhWIC+rL+hE8EweDGGgqsUT
ltnNvl69sezwdON8zllpGHigURONqaAW5BBmHM/NHpLzr5Sy2y0AzKZrVOhXE8k3DA601SSMFKQ/
s6yjZe/bU5tAXiDSbAUHLhJR0Fsy78khGz6kUuBDpF5wDACdu+iC2+XkIky2Yd0ikPPPCoiL/ILQ
FEg+H1xmAkLurDWb/0NcGM0A2GLMa3qQZ7UHh4DvLJJTMWrHtmd0f45vj4wqPv3WZkSoPfm0x+30
5AUtOItSrCdRAY2AyZNMlrBxw/PZePJ62KnyhGEdehiix392XUqvqh5J7NGIuETVJ9pvdpJi8rU+
4hWOdCDsA3NGlC9IDnJvRxb8FAK1v1CjIh0RbvL8Pz++AwfM8P38zZU6y18FtQLpzwLqlvjMaEGM
U5qYQfTDawJJ+HuOvXUN7gO4FZDwhFCDaqYt7oZ9bZZety0Nk1841OeUgv3tH4VDaoS/xWVdODT2
yVcx6KbZ/vXS6mNFOZgzwIm02mgOVVGVlRma6JShoo+re5yv8B7OxuEyphNUUaBqQ+4oLnFHAIqV
65fTPKOETPrQ4rVkThrqNwAfn2oGqi8XH9gLxPTIb0bP8/DAtoURYfcBCdh/ZMuVysd4fgc14jjx
YmsVlRa/nMsWa+fQBBcAd9LIW7ah+MLB+SaxqbZ9HsARfFlCrPWDOWJ8fk0FNAw4XhZMe3iwURbb
BeE3/+FaB9hoIPQTdTxxZf83hFgOzktkeVCPekbbaqsX90jWhil8SJgi0H9OX9uBnyxqvt9EuSZR
xA3KPttQc4ZDgDhK35T9Y8uLzIjgdaP1FKn/x3flH/rbe/N08CMF6MXK1djr13uz+iSF0anq4heE
zu4IiM+U8ACDuCLksri2577lHlYXfUD7PLREhu2TAW7DHtqc2rrXJWFdAUYIPszQQeIuXWKlfDlY
U24bMzrswR5Jh7V7JdMnB2RWgYCO2YxWKgLY21VqzWD4ZNGAbRuRX7Qig1rsgCwR6OuZbZY4JwE5
GzyVn47eH5JEkas7N96bDo6JrQBQUM9ZLVCw0JIho5WNlEROpZi9h7Fe2V78dzWnaIr9suDUQ6GH
gmNfH3mp5P496Vvoau31B4Ciwy+TtdLKBF6J6oCLDEGLxJQurPdSb/6vd16v3HRx1kbEENbDL6sG
qPcpYAKx3HAlICFE1HQUTIbyr311lt0cbXYTSQdwWg1G8nitV1rEG/XiqDnmjwNi9J9R8OjnpvwL
XBMNE3ELpABzcBfMhte1Y65Y9FY9GcktID1AN1vTBwI0IM7TMhuQHw3Gh1+Eowh++v//jafsq3zN
EaEsL3omXIqVWSD16dS6sJ9WjAYAZLb4o9zOiFosMlKRHp2MSMIKaLiEaz9GaPKaNEAqN8FZpTyn
mdDUZ3KE87iMQ4ujFmwKRAlhnanH9iYJ1QVYPT6g8ImpWpSauxCquHqvrXj1mN2lc8Ojh4djsnL+
Op2cubtEs9l8cwgbAjeARqgBkLPS5LRbYjZZpapz72LI3mqFI7JH7oR1WZVPIkvi+gtUemInu7UH
toMDDZZgpjvHajfJoyPYoPqofyLww+4FJLGqmYYIb56ICP+3SVdh0/qEtxQAWMkMT5ggtnsMy7ZC
0cDAbBBR6FtGWSAeiDW70CcvWVkwyfNsk0uNwe/ELoaWAqtR91r+5LLjB0GlIJ0zWB3/RS9gn/X2
00Q5xePzFzY41M+CyYIdZBL/nUgxNPsZ1gavbob5QMevADUVVka/6bf7+n89cX90RgyPK4Jd0adS
eRkqao8G5DwO3Cftt16EtdhahvnCfJ36EQ3w54mE6xiUgh9S5i1YB+jgo6cazJ/A5E4nR1g24ian
SzaUyi7OmJ7BKdl9MT7NF8apj/F8PxPAXegBx/DpGaoTpDRq4tHhWbEFdj79wgCDy4aM7mZPS/Cd
vlsDaNCwrer3wnkGlsYW8i6X1dV050knpnoUwWbK8bWGDbWszh3DYjeoWH2JLXUvUkf/acqMD/9Y
5CSRLSN8qIBmaP7Wnpy/waROgH9ejqJjm5OuIM2deUXKXbJXAqGs7F32dcVuigreAGRAdJCx0QEK
MHzpaBDQHiN0r5AivBv5Hxv7Fjf9lWMKvYUFr60XVB+3O99nQdj0znCyxLGVSkk7xY3EE3tMV55X
pCAF61sPbaPcg07mAP0IvimQjUTyvsnuaMkmioviFNWeusQvNbgvr8afKqaG+1meCnU1Saxr7F6U
avMdpHoCodulJRmLLcVfIVzAI/IQxrFTLR+uKN936keI/Zg9d+j7Hm7+LS77cU6pyfTlkl85x/jB
s/7L8VofCnVVzPaaiw4uZMzdoYNxxcgn7noJS3i0PzlB/R4Y6Vsfu9Sqsbn4X8STzr6J9J+k4hz3
mEhtdgG7d7h6T7/ljUZwJ7zx4K89IeUTeCx9g9YE790EAHR3kW/1R8yfAy89gAMHnRsua0hSOc/u
VCppowEUr0HUYTfBfrzVz8UvSShAlKBmqoKzgjbz5B3csJbzDEMhHJB7sM1H1e+gynPBG8mRdC1l
Ywvzv4sRkrJvLANA7Dp08KkW8wUVR25QpmEk9nnaK+UYpWzRKwllPyRe5CsFBdQm/wBxL25GlsjT
ISrMGcXUdlFWeZSsaN4Zpo6oyAu8hHnk5TmAVljjer4O/f97L7MRBqIlkR7fxULoU4psltd5fShX
eoGwWW8tbY4J+pbSZMzWJF4jUcClHFbvEvECw/ooFU3wQ8wuCJvC8wfrf94gnYng4fTEzckXyehU
VXB9CMvGhr5tWFmrgDW4vDkVvpihmWsSk3U1sjBDA7upeDCR1pi8GtVTMwLjO7b6M4QjJrPNCzn5
rkbC0CKXL9sfuTfS6+cIciD3CZ27X9Et94v+1Gg98T9/Mc5yOVZOgC8Ec75td45XLSYWSKZfXm+M
0prYWs9Uv8WbdqFQbTDM9EoZAojY8GchXM5W4gTODUf3uonyRZQqWhzuqzTJkWDVDD8WKngBeApD
VE5FrBsEUcbPCOBGF32v5pR7Wq1HlaXAA8sN8bElJX8uv8u9/fBxWf5XJmBC0QkRDacio9RVa5VV
TJQftvTgAIz2lFDPRTMNl4j6ShYUBZ7KsR0mSAm3BAXTK9+MObMS/7CW4HUg/r4SNX9SbYkUX6Yr
4pYLFqtOcwKqvPTP9wiLrFE/lSclAniE4tYdk1MqrRI8vTBhbR4U5XC1NvbfZIGbCURPxdzOJcDm
KKqrTUkaBvE9RDSoAnNRNp4GEqtT82mwPCpj9fKgYIMN9FD900PR1vuWif7zQOl8uPgsZAM6wFNp
I7KxidVFlP469WWSIli3PUaz1snQ/F19cu2r6htFc0b06pdsMpVN5EzNpaFnsaK4GAJlHZQXjgB6
1kiZZo4Yuv3fQzeeDT7Qf7Y6iaxb3Y80ktuilCup6Fb+s843P4RlvBW2Vwrq/dEhbnixKy+dEPEG
AzApuBwD6pN4VzQttdhbSKZy2voJtcD1TLsGqRwOXagOPlInomZ25lMg7GHK/6WmsYoa4lM4sml/
FCwRiYfeTDK4NRceY6q+jpUeGZ6XZvO+7YWGBOfndUJZN8MpE5T3zqjr+mpUubM38xzWeoPw8ayD
XM6hgRHnc0RH7J8IQNB1Qtr3ASvGkVrjPgJlbx8Sa9rVgYU4fM15a08ByX7ddOr5UFUgiOMw0SgZ
zWBLifCChj3t9OYebpO3wR7wt3muZiVABr4wh4mx2TL6kb1hexO6duuux4fzXnNKBV3oPFPvj/n4
6uJz/ECy5O79VsMG/oiKsEeGPqhj6BeHnLdT3lIBm+590mQ0PlGjBeCo0G1rut/NXlu1lU9aqFsw
pZJwuPd0y6YuHlAV4fDhC1W55281C5SI0Kyc4gbuU+V21HAjqAnNtGVbjaghOqgICflqqhkKEmi4
gOmEzOXRj2bOC/rDPvQMbW0aMF/9j9Q33NptojFmWE7oVNhR5nFHgaUXHuXcaPksI6DlfLAh67sj
IS3+VxAw6AWRgWEqKbodIguq0Sy1wHL2izXYPLgs4VkjXQU9dnuNbId5BPMwxNk/MgKPYHc7FT5Q
WVqzg+Mpejnero3z/volB0vY/kRQKyvj1GHQGJsO9S1YuDjYQLyKsoTZBJCSqg+7o8fE2f0alzLF
sUv0/GiddzoEJrrimyNaHhjDWdtScuOY4ILS1bxs5PZjQvXE5EF3WAHsUNIo+FdEmBBR1D7Xr81b
yz6Wimt70sFiHxIeiiqELKs+DYqzFTlRsEJ/Y7PmK1jYz22IIvnibVf+/xIjUtbvlIuzfmyd8sHb
VHoxQrsTNhyF9JdRMgf93hMwzBcxCBl1+I+SrFXJIqSX3murXQ/OrRa6vyWwvwcBaxQwDOX1smcu
MWrMMc0eX4gD1bEzFyPOikLSWkpx1e12yHkKUDesLsiRPQZmiD7Q3GUN1FNntwICHi5eFqfOx+ng
aR1SvMHGN4FDZnV3duc5vjCrt9z/O5S+Nn+kmYEWiWOdC6GcpkJbDGGL9OuJY++QEEDeEpg3iVCf
TueMiLe0ls16bfvPp6gNmBC23EIpcBf3A/1guzxsFNhFljip3wgL/hl3SuwkbalodaSuKUxonsrK
QJ+jpGraJRGCUG1E4XBfNu1r7uePskLE7IgWUTU9IlmvMzPLinLBHTLevdgUM2xIuJ7EVP3jj1q7
3UJ99sVFHPRvpBoEgFU5QY4OUFxBLs5B/mhliGgoiMEb/+rhRVxY87mAGTKvIiCusj+sM3AALeK/
v72pY0DBG1J0bLtjK2IODnwTI5qdnZOrV/7j36V98LgC82X+67L1a4oVtfG9VH1vJJUkFac9szZs
RVZzQZoB9ECqsUExAXCEx0CRENqnYfQrogHBLgkGXYh+25Ub139uQJsHlekkT4BAbKkXvNMGD2vh
wb7srInz++jNdHQAQr9XDZNbkcGf2u98+6eXQwcJ1F6JfCtyDU5AlFcOIfx3QDDVPT8rtpahd/Ej
XpsUCmnnj22iJcAqQqJdnaTcTfIwr7M/4I8Tvx4QdCogm2GKsVgK6vQ7RtuAKtX+5zTDpx+jVY3a
TRKNXDmdgTbtzbJvL4u0rB2DSm1AsP24OnbeFXdZ8C1gw83LknvCEQBA1GBxPhOcYsphAFcHBL+p
I4stdgdDtiCjxN2CE68mbUn7PRjMRk23f0T32SCjVHXkWVHnK9DEr+GRIFwVPCktCEOfi+KqS9Nw
P9sTyN5SnvJTUuvkvQmVSviyQM1TvY4FdsmSDqQbm7eLXyF4PAsJyjSPdLuDKVx1J6LG5Nf5s8fr
fIVoqONuJfP809VY8obpJqXaIvm06w1QTJJwKZuGz3jffYTxZDZp0Z7SbrP05zzihZ89oDOLMZTv
xb1JtFXtLqFoy3HVLxWiV6ZE0M4pEPypcaP01rBZgKvelV7H/uK7GjnXRF95WLoBYcxRFbvNFXFl
LyBtz53rPoeD/ogNPGrIbFLiulYZIeMMSQyAXpqbAswFuu5BXIpaMePI8wSBZwKLqxJuu1IL6Mbj
rn7IuouHMEF2eb9R73MfmjZ7xBPowkROpXHIuP/1jnWasH5/a/DPZO+lLcNfC4fwEAbJPZmU6eIE
eOKR21AR8Et7LAbNWL+AiNLbcFxF6WzI1LueKI06ykbyOl9ilFD3eZIPfsuflBkgdbP4wlUnlrhK
ECQazC/qNzPTq6F9skPcq0bmAoHVgRTK6sXPTYLDABrAgt7Z2gVeGAxUAHLsnzo+6r/kbBFCpAB0
+7XYWSqOhusmZrlyMiyPh7AeOjXIsJiSX1SuWaPOTyVzxdqcmzdoemAS6uW/lto7l1t2vyJzKlm/
i054eQrVcskIXmYKcGSjskMWIqn85xzsfglCWMoqu/qGe+ShRyoHe5b448ctbz7UzSfB8EBe8l5c
GtDg0gE7O+WwAH6QbUe4LRwLna3iQ2m7FMA5ukmDUsONk7zIZQuPKcq2iTcAsE1U4kLRXNtJr0Ly
PVDXxfPlRkrv8Mg9fmKL4Slabsr7c6F3gIJcPmvxcsOPmyk3OpRzmVpVOiHhwhZH81WDBu525CxV
OfvSzxnQzSVprqL6NrXIhSHWO+dIpByA50vyKOWnGraObUU3Cg9VDUkQHWevkA1tCyPI2mvQiJoq
g+mPIhCtMAWyXirDjUzXpm3X9OzcrcSmhMWlvM8gsDWsBOwYGLkqZRt1vEnyusuYXCgEReJlS159
1+/K8N2guqt6C5B8ZRaFPdoPcrd3H9dPCHQzhb53Wx/cPZ/YuIDj9Ykp9WwSCWVmlpV0vx7hPm8Z
MmS5DVTUgF+PV4bJKKYrpRdSOZZPqeqUDoW1yycG9LsnHQ1nk2FxmJt9Lp9RT4BAUGe9RZ5RdnrO
OeVjfDcrDtMb7eumwCCzNjqONzwFsFPoLqHi+P2Cn8VRUjKCNInuPQlgAPJKLfoNFO4mBd1Db4J+
Q0L1U15ekqSIOVLPn7u0B8oRUmxmCcR8Y3ZiSN9PB0IVO+m+Qi/P33WI8P5yPxkMK5BuJIqbd4L9
TVS7QOhhaA394Rg+FzatMqfLiFipqm0IrA1ekKYgHa2K4z8ESKY+Ng1XYkWz/QPx1FEKbBRNOFXO
SGB7N+4NHTdJokz5qLbJWql4aU6oc4dnImy+8+zKIM+iQBm06PYpNUB4qjTGPPg/yLNqHMWOR6WB
CXz9yPVFtq15Nobg5StOM1zr5MFSEOjVxFgI130UPvrsYUmjvr3j5bnmwLBzlo8ptNj8FnYCifRS
ZXWWv+X2sp0GwXkgZjuDloIUXJEN/lGhDpGheBoOU6fkNGSeIiV3eLESD5Tr0W9A8TLAHg3lSo6h
z9KD7hadVRPIhs/J2snIa66G3WOPQSDltol17PoLOassiec/8yBYttD8cRDCxmJVthIyELRkBKaP
ZBjqn8kBWUFCkAbQvr2zu0P5XEg+y/nQwf3M5D9FYWd5O1tZuSeR7s1bK8tNQu75aKh+2dDHF9K7
CixM5a6WMWGnFtUP45+aq8XWRtzQ+REtqb975rlZXTbbpQMVjqhPXg7mQH0r8ZE5/FbvhQdmGpLE
3sUhHIrFDdcpVHrAsXaLSSM8PqtGC3uWf3ztuzrNydRE3gnjWoJ15HxI7ENXSOxITiAKLwc9VcWU
fRcW2QI7hZ37xvKkjK6KlfQ31kLPtowYIQx+qiYtytsNndK0TuPrZpeyEOMFN4oyyjZtrtO0D1km
p2Ju/MAckxHaj6X0pVOwMwrxUb4xokCJTY2bTzRgrScqzBpTo0ZkeV+wDkTbZQ7l8gNKeH+pfWOz
ksuC96Y8RqBFgiYqumZBm3D5dYeuSuB9yOAKQv6EWsFIVYMGypgfNFjaMIT0cOWUm2cA44bE4M95
LHI6FVHxRX5hk/4XR/M806Vj8WVIwoDqtg9IndV8HbBRl3BxGUA/clE3yCqRGuKNxbf80WiRtrV6
n465ANX2nV/ltsEDuh/NyVGx0gAwI6gHa6Ha/IBuI4Zpssp8C3iX3fXrg9SO9HAztXV40AjJ+S7R
O5GpQ7KCVz4U46zhQNeFveipaMYXZ9GhpjCCIqdUtSua4keXGcnb9aEXH89vrdYFAoYaBHOSpq/d
T3Uu0G+/B5B5AjtBakhY4HB4oJ1X8OSqVA98/mYhOlo1419ZqeINUR00e+pY8ndCoObo3IJlvclX
FW62Q46pn1+u9KGae8QepOMuuAdlvLqq/I3y8B8e0CAk8zatxicnTHyRgexNVYwVI5SgRrL1cc4Y
U8CoWSuMtcf58nsMCOhTLCmrhX0HCXrEtVuEl3AMO3giYQq6bvhXUz7J9EHvZqnl+Xsqzd//hjvE
yBHVri5G+At0gGva8bN9HDMRdK5+kPFaCz0b7yHGH601L6byVLMrZQ7Vxa0LdZ2rdHTrrNBV42Oq
/vuOmIOC4oKs1Z+0SS8v76OAg75O8ilblsnTa+9EWWkzZm+NYuLicSEmsVR5wiQiO/x1zdQoc7RP
4X5JAo3wpfFwT8TYn4ZhqyEI6KKryiSivyZwR+iZt3HO6IjWFwTuoGT69P3DZTbAD4GEv5QDcyhI
gxER9pMhNgMDbAdLaH4XgWSHOsCX+ud4GOBsB/gbkIvxFHDkvXpvA+GqWiJKVLsddR5zVvGyXfCl
1SzesAkOzgdIY0LSB08Kc0eV/NMV274EHIH363kotCyv5BtDuvDuJnWbSlXNnniODXx10D4loLEf
c8xY6q3W4GJ9oW3XRTVZJk0GDbTvFFGZjWk8B0Z8e1wNR51Ar1MU3uY1EYiS6AIpLmgmy5f0ZxvB
eGLvlyp1WF8RalIgL0Ld2q5I4JTFnBR0s4XO2uw+xXuYZthbzYPqhTGVdVhp3j8tFvwcouMEnR79
1SIXwjpiGf/eTgCPkcUi1EIIXEBYW4iVeQTG/G2fmpzwaDSJ/DxhxqClH0hmM0/gSLqgOh2QibP1
/1sxTLDYDmL5puJxfed2s1qpeSbJJcFEvaGAzaafP0J2p6dJnhTmOfkDwgbf+jnLGS7JMWLBgIUn
R+vKLZxPCX52Ij7yrSfi3OTlhWeJNEv4ELMBVOhex1uCvcX/tCEuQXTtuPWm+0v4xv9RmDAFh03T
vBGz9nzI1isN38b32iz04K2a/0WHF//YzAdZGTEAwCpOYxM2Rf605uYfHgDeCvFJiuW7VmesXQtd
co+ILLMls8k3Zd9pXq8uaiq5D6RZW6hAZQqhd6YBiNpRgmG4wgs47P5BEm4HG6UQ7OSkURZsadW8
sbZInZ2h1zIAj/qmLAk8HI4oijVTa/9zHJRdrewGGkzqnFTYw6LmtsWPUfg5QnIGAoZd8GUeFnBM
aSJxIy2JeevX4V7knZxtyuA4O0sppOAzhJCOUIRvjr6Ox5N4ORxsuBgGbgXeXZHdM797Ren4JIfk
OJ1lcH//9k2i4TmoHX9D9+Jkdt5prPkFMeC/RHx3XidHsHBs8pGudrFIgR4x+bmfI4ilHq06S11C
ZodNSgz7jdimUEm68I2jrtnssDCeECYmrFOoWdAGDdsr8mhO8/p3cIlJUCxKuhfv68sf+sxma+hj
L6NUSKlARGMhxYZGUJ2hFg7mlaS57DPcBVqNHLNno648hDGB0k6GfMnbA5AHXm7A4nUCHFHp2D4x
2aJtOceg7DoDehuvtoYb2NRiXPBR5UXAJjOz+x3Eegkn6Ux+ORV4GVIsoA9IycK+ejqz8624rP5t
S3Jg8J0r0W193f7rQ40LSotzrkKBVbXxMXMNSroJ3YDZWeIkpQMpmM2U7WGr/v/5wUtazuOUCv2+
x6ufP5TDPMczv46k0rIcWM+fNGpeHoFF+36Ka2CBlpsxgqh3Xuryvgv8n8H6YcDAwea01KtLy43x
v8CWmWcw+rGclTlTtanCTkk/U6W8RG7hdWMGgNkeVc3YapSzrjq1KDYrWEq5f6/LxOQnXkNL7xq9
Cz+e95BbzO017yUKMJk5ObH90huacXZDldvNiyXHxmptqmKH6ZZirZtHxNDfPyYBK8aexe2cUzcq
7/HEMsBXndf/yzgirshN/uK/pbf9VvPAKpsS3rBa5HzHzzCPpbzPBGMIn1mBrwNtXUhOBPan66Fq
Sxpl2WwnBypcBtJsCaqMDtYdiqvE1PyjKIsGyIOVaQJBbLTOeLkrefF9N5TUjWytwLuE4Pp0Ddb0
hGKefdnIJ6tXJ8BlLLwXjbtdB4VKRGCI28SlEjphFjdfgJ9q2WJsMQ8ICNUPZPAesYX3XGVI2FFM
6cRVugcNmszX7HP9ktrftU67Or7A24bevHN9i1/NQk9iB5JKtFGiVEuyGrFTDBfVo6Ynix0L0knm
dT5dQprJZwPGPor+5q15kcwJ+qvgenaV5/qo2S6qP/9i0Mxy8juOqL16w4+5GUetgPUaVZbnr6gv
a2y0qHpnqq6cBmip1pg6H7U87jng0uGXR2PUN4LSLItRXXhysekySuoiZLZFECYRyA6hVfYXeZyp
zf4gOlHV8Z2qmsWkTNORU6bOIhFDZCKQDOhb8VBddsGKffuyAKVzoGKSE/vITUIA2ZvwUNSSjPxC
8EWBgrwTUm8n7CA21mVDvVJYYN/pVhWUcboubFCyiyZuSnXwOmDtjur72AsiVPI1enRfVUIRldiQ
kqdPhY65OTSyDUMkHZiAqMBb0aQWYNqem2uv9fGrUi7i/UOF+T+eEisPs3SFstqFijLWAsbNLCfP
4M2GvjL3hr8jFpmSeQwiATLQtffOPzS+XVFbn9ID6F97+w4tSDQudDTMgwQjMxdozd+or9zM0A/1
vsfLMX5z6POsiagEZ54pdVHYF2ZcPKJruIv091z+mjwAtQi2jk5LsoRS6kB/V/i473L+2fOCbN4L
Hzskyh2yR1ah/1aWG/cU9H+8l/2C5sen5iKc7tOZ1WUpBgnJctqgwRoYSFg08lgSga1WviT/MbZH
LC0t4pkzEYmiHdT6+sYv3veL8moS9DMAMkrlgnr1WIknnk6J5c6jR9YHqcTHsOIwYy9VPywvJilD
AAyyGnTXL7D+q59rypmK9/gKpjvEMxe1G2TQWsnAfiCnVKxcExwniaoLRolY+o7vLvAhjCN1N9DG
nQ5t1V3ifzY8j3HIOxIzZuLNhNuHgKEwroGvjZSN37kppHmjr0Y3BinrG+yuPzyHQtqN/j9Lzx1J
+6/ygIfGLS3kJn0ijeqeGLyov3uQWyEDduDBfo8GoB1n0rM9A4452kqdb2Mq8r8DdvNj0mdBygKh
24v2sLDWC0w37hmNfk0urkD5XdEuTHVmQjx6nuMzhU+3uSgB0Lgdo/5lDWEnAhf7AVAf1cH643CV
80t1HBRR943vJ51ykILMiFFaQ/PF7L+qmV+ePGaH+VyjK/K14d3MZnsqiPdFTUskmP4Cd/YzkAz8
PX31rhTHAKxFusaxQk2F1Q8gw9G/cmCL738LfmXp/7lQEW3l1vmzlaE9/606Iv//9bxquj6SpgQW
7UNng+xVd/thfHM/q/pWY8ahFtfi5lED8TW76IrYFIpBMMNrHVbamgDf/YBMHxl0CjffNY+q6qnI
cT68xR00hVypA23sgoNLzvmIvKYvCxrqZL3WsNbxFFJwazUROU43shsZnCdmSqb8rApNQ2G1y7nv
pQi0t6HWnpo8SpvymFpbosaRyHXz2oTzrtzveTiLcE8Zx9l06DAnsA8OX9MbTprubbcM8iIrndkV
WAuIzc4IUIN1YJhEkqx9SGKpB+uZjXu/a15B95zMJJmyBhHbtpcaUxKgHqaNbGImYzHuzJaW6I2a
T/ioh47uKoi0+SwSrZQpfsYSVfahTwfTgsVHvbZRS4kkI8jh8PRi1062UI8rwPtCzFryy9DAo0Sv
5Pw7qXtmCCHzsjp3UvgFp2zqpQ4+rRTV9wnY0lxstkYSeNuHwRZgoCnY05LSDJtmFvod6a/xVZSO
uwG+lC+1ISfzKFokrNanMqKI1SpU7TDLkHOHkHudGCfZUW8kpS74qOKuzxq7+Jxb3SSivSYE4D0A
DVxw8dH1IpeTN5oEcpOUTvcy/YCDVS913fy1gvElgOSRGX7F4VsovW/O5PamY6GlcVoHfi0eWhUO
DaK4udKTWlrF/x4AJpd3+nGKgCZ7lZm+mzStT9NVzFOkgo9z5C0NikUJPQwkd892ChnzVRdbpD5Y
q+kXUTHxupWzeMU+3be1vFsGCKfEj9uhAWQpNZ8FU1bXZlgCmSZ8vb2C5dvd59JPTckQlk44lyi2
3jfGIK6866nASV5X6550FHGh735HIIBIkncJaxivFSLPlio0ElaDyYpIyREt9dgVGIitMcO8wyQj
zBIH0DzngbdndNM5SuxAMEyYRDpt4vImiP36M2L+9RiLOb+OMJ4GHRqsasbFOLvbU4hIG5GxKOo2
cgIhG/oh0RKI5XI4rAzZ6wkUlZPRFiBWAWkK7g1tIZZZeRsdmZT+l6omEl5UbB422sz5L4O6kMRs
QF6FidXCRXbiu8TSrAdQhtA0pJWdX/oZ+KiSlXTQWdyA8/EoOsb7sdXW4cx8T9boRVhNXn4/kUHv
54q/yEKYsk3TSsi4BTEJDtTAM2jPPThic/aHex39NlIIMSdt+3bK/SC3fN9lnhFAG9a6W67vLX7u
i+Xx3qW6uEU25n5ep7zLjp3nbwrt07CnkY6pC6SKOBAZv9myO4yg7xIQQwpdxVjPwro4EH88Mr86
zbQR4vsVLMV6zFeikh+37rrIGE8zt3VLz3sKxvJU1Bgpp96XLVNsaFrW4hQprwEwg8NIRyPMT2HS
lyISVrv4a2Vp/CNUGrEc8uQkOMRgWOjSxjaex9UvjDMCt5zyOkzJ0StZQ/aITzCj1tv0YP0YDJTw
pquY/IIT1CkQSTWnHJ4lnmcG4Wq/djtxYIHvB7o+ZHue7FP4jVflk4I2JgdXTGGN9x6rpECX6tRD
4Cvwam4lJpadxcRWCmjB7ZmvITvBuUXT8urJonJHC3Pd1b37ET/gfaG1GMcmynk7lkkyDt0vvqP0
PjN1zVFEPzXS98B1714tz1I2OKeDPt240TDAXunhuzocdjOzInkVOC+ThHOey5NYm5P/IoxX8y6p
uqGR/Ea0i6QHKPEtF5UKPZ63ibmRgdYGWmNwZX+iDL7+4Za86zyJ9G5JyVKQhNnZ66FrcOmThoM4
8yL5XeFi809Aevw/gEgmcHULeyOdz3DpMdMD+EWby09KUVurCcRpkqC3Z8Wf1iZxW3hDu4wBZhbn
c/pUVNNOvnXpGUjDwguZltoErO3YWpedfuQSSBSU040E8h+eG0gclasHK0C7J9y4ClX0dM9Xkwfn
wxExY83CxWMEgnP4MDBh6WRhEUWudg9zL4vbAS2yZfJn4E0lzsR6nQvfOF1/69Fad4Vimlvt53Nh
fZvI9H6rq2t4yfV06mspVcvVMks+7ksnzjY+d+jBSMwRvl7MWpXtHkFWUBPm0UP0P2GtHgH7MVwL
dGyaxHjcEgGF2PL97RnTcHx/U5fgzhYN0wwwel3EOj9dFXM/y+GZclm0NfQ8J5gil0g2qdv3CeaJ
GMUkRf9upJgUXgVh8utKq+Ce2rxFmFS1shAxhPUfoeL2zBgZqzupR7CiY7K826pBFexVJENUaZ1O
ahU6/U56n9gMxjoeiVHttOjnBLRdap17ZpMPgWOtUdEdGdEDhEdhibB8v5lLmJBAZ+dLCOmVP9mL
4U3NhRLfGk0vMTGzaJuvb8+X7FYA+V8cXYlDZZez1FJcj3PFwcu3QInd3OsORsTNZcvBpN3PYiH5
Vff26dnAhAIa1XXB4mPW8+YjJepMUpeYWcXVT3zmGpJw3XPwc5Tj/4zq7HI/iIQ8cCHjGs4dV0XW
oo+P6Wj9pU6xa+tU5fmNL8fnnfCWS0j+NHs8goWH4qmswOIOInsdKGv4XFGKfzl5C71SRnYnDsH/
uwioOYPyJ6m+l8jT9ozaoSVA74wvJLiBxg13XRFY8NM/FfyLRkcKrrE3Lf9k3Aegxk1VYarlLrO/
Kj9xIQBt23czuG5cMDyYcBXT9RPlKQL/r3tq9hjd8DOA0fl5nszEADseIJLQNNwgLpJHhlYO9CoD
w4tyUqKeNfOGIHM3AMk+9/Vrxlg5q+EuL/6RsAoNmQYVTiUyMywGloK04pxxhxkm+h+1jbbXsPiL
Clc4SR/Hh4PxiooPE9Y9YAkbUxL9qK9W5lVG585CG1j8f8EhPnXTj4mvfYMwCHvyH6xO6c7FKbEV
Yo/1ido8CPlupJ5op4KJJDXzb6VBTAisSCGIkbV4jh88Ab4c/bsQ9AK9hwBWqcgVEAgrdNYAsJp/
6dXQOvzXjQGhJb1tcmv5cwdftQB9hCvYcEi4OTHNGsBRTHADAbq+R+Jr+biCPfOxNSLqmR5BAqGN
ks3cytcneeVp/3TBnL8x6pRx0vCh4ZLqecKRMRxs3zMVuTttmUioWSv9dws5Cslvstt2bHi55mWF
gc8xblwXJcWJLIbew1QkcDFT03hgBvQyL7alB5e135WgvAi50K5PABuVrSZjiQyzwwx5dJgIDPqd
iqfds0teTYuZnZX4dg8Kuwf446X46NWvOCL8NuS1R4cp31LHp7TwaIDfZHLDHmZsUQzvExL6vJNz
h7CHG80Ory0NC8M7gePmCX1WG+alMQ2X4Mt0qA9fdy0uhd8XcAUOfAzG4zsNvb8MtmNAqyUGjjK8
ilkVuHhwpISlYcHNt9k4UsDp5hVgJ2QbbK83YxcsVv9enhgmyr+FldM08S6jXfu+81BUC7c0/FV0
85MWjoPL6WfLTqzfKixqrjy2JE63/gYQguNSzS21gQomftRBy1bw2qtPJcdO2iXGNHitXyhDGSUJ
0LGF/fXvTDsVKKDsmKxkvtsDsJPdA9Oz9esHJnPnhmoubM3GjrDvQslsQQJ1LtIHVa1oXeA3mukZ
awrnW6ur4OJ5saWFrg4dAOeHHwyzDUmPH17fsP8vFnpk5ReClYw41FUoPl+YRtfheSWupsjzfjEj
REj3v8+5Bik6o2g7NcGnN5GQ8nLHDr8hvMroMwvejAFXrfzN1bWgV8WKCnEEqk4VvYgGAUhvpHup
qT/ZdchUr98nt1GvwSdpNgNLw2RIxRa0w07i7YHmBD+AgaZ1o6+LX/cBARlzdQJosQJxJnt11vNQ
WtTxNBXuTwg7SoCSWdAPfvaW/nePSCRkQESkW1BEUXWz9eS/3zSWp1RwLn17jkaBuOW1pIehpgGG
mXUzGH9mH2O1OVnr4tnYjW+RBDNGgfnx2qvfCM/N95dr7NKEoX6nsG7ZApGlJ+DKFSC/U5PVTuXo
27DgkHwG/mFfuvFB5yPRrDm6CAJaVSnkSbz7Iv5GfB8cQZJK97sA+FXSgkE0MWBr3s1jIe1F/VtL
je2U5fq/h230fP3AXI2ZLnZdXCyZA9dFF29rb5X+0kqW8ssLdDPnUoPOhB6xAVRnDl072F17bDcN
/A9ULj2Ry+jPdfvu/6EUttifSIYd8d8b0d0WO7uZaFRGclbXU7wg/cNQEd8eQfGrUR+eCP+DYC8q
m12BSr1IeuSsYsvONhcKafk0DWYQNUZoTfFaS1Y9y2YOjfX6jggDdTq1HjZzxhrE0or5gmUsMlMq
3jCCC1p5/82ZsWej3HskCP0riXqqJUStN1aaTxWdXAvuiGRrebRquW8XFtdecIe4di7bd8agoHos
yJSZgiWt8lAlP2rERs5S5aGQr5PNEqgppdYSSacrlqREjIWn0xZwDUfb+hwkZ6VFJvVvttJNtJFu
fgmvvdnFJGctnC3g/qosrBXtzoHqRRavC/kaw2HJ+uFkj4T45eO2JKfQf1M1u/OhMiaW2hPeppzk
Y9lqUSw9gqGYXJbj9cZEVX7zFCuviQZfyXXnWGjZpWPEUQYZo9BTJYGlemDfsxF1b285JT8i8rFW
l57ucNMnOwAtYMcKUmNuidYs0iislmemMTJdxtK0xhC7XZWE4pWqdFqfH57sK8CDyRlcEtH67HGJ
90QMAy6JnCjuFVgRnlaAnAMMHckbjdeK+0oovdwKundLIer3yYlB6KMLbrPHzLAVNCt22kJO1u0C
NravdgNZKLXhDaVM+nZ2U0DNXcN3mf9WBu+G9y5MwV8OjOgU8aT+uIsnt7+94dDuavjEopvwhZPE
X6d1iA//CQj+NDOlmGSGG70o+/5kFbfskw2Rg0ExJKgnD8kFQy2IL4dFwLCTdoCDxSFPnVvTiEo8
wpxHYjHdIr9cttOnhNpQ8jLyKN/gcxep+DFnfxoahjG4aWjSUxRP3V+I+jHweWc6lAQvU99B+cxp
ndnDA3fz5fC18gIhDAht4XKCEFu8NMMsgxqBLy71JBg4CO1KFUB6oIoFrrto2Azf+OQSop7RwgUM
dgIPE/O3ZyMkuk2r86BpTDkbOI9Wv6VEiYoTR9lQChd7L9qbDkHZt/9+9lA7qck8zHjjfgJPZ/KA
juN4TSQQdOGbVQ+irelz2wVEfL7b8SpmA3CBBP7yKFPwWEX5U9SATLUcdj08OIiNamE4jLCYmG/T
FVnLVWWK+5BX3lJku/jDhlke4tvglZdTrIXjkdWS9l60JMa6Xatf/qol9B8NgFnahFqY+wKh1OKJ
bOMoS145KNJfHS9ZhWbJitpQwHW6bijIAQjrbUIGMWWQ97mYsyqwQPsP4VPyxK4zJsEMkKRAkEG7
9u3ILEVdvHCU7vmP7WGfkc0w+aP+Fxi3Upnx/UywceAlcJZG6UcvSKVWlQpgnE+JATFPGlWnpfsx
a3Dm8UwUXoKcXaG1T44ixAfLVTlv1RGqYRipdEh6NU89S/HSoZzQQeyNvlN6hU3Tkf7y/HLffgcQ
JqwKI6LP
`pragma protect end_protected
