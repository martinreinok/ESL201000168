// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 03:52:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VEgqp3Un84Ii/2vuMQxfDDPc39/FQOPABpkM11auyRu2QQHFbUEAJPXY2fSvEauN
80O0GOl6U+7nJCvSpxksvgB25QcLFT9+xvWLJcITnOKEJsSaHGzfmKToFfWaeKdy
PO23jUamMacF/covCcGA/BuO6QmZjNGbNpkJ5oIgNjc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21280)
xvSsX50yqmqsbNI6ckZTsjWyaT549ToIuoLpmQ7fXY7ek7NtjklU7dkV0deO/B3i
Y7gQ30Lyejgv7Faa6whbePNDRxdR3o8WQ18uDiHdsThBAnaGO9Owx9sSa9lswQac
IxDUv3r+rHUgQarzuhw+U+wmtIaDS2LNVcQJejgJ8+cyAzPLw1EElTlaKXwojAyh
3afDHAQfgdxq8g6eyOran+ugkZEXuCL2pwv0M6kl5bj5y+JS9v8naiNFFMI3/OYD
xNoFy+SfPyL530JJTCIa5j7JQnhiQ1Y+9sJoQIDhjtZJQKKHROnanyp67K8EHEY7
TYF9UHJtoQme1yPBNjqW0dj14+nwX3jglWuJSijHrVrRfhMHtqtYsk1MqPPzoCCv
qyg8x2DX1+DP14L1G4sPxF45mp5JX4uS0X9If7vV7mE8ZTe/uaueZL95v2SuDgNQ
OWhmiYMsWy6NbKsVFWTOkD86T7xGkq7xEa294eh/LdQkZ4jcgzTsSBhM1kBd9NfD
7ERcR77jFL8/bDm3r9j2vK9pAZgT6FKRacIEA2OGkECrxzQh1z23KSafQL8baR8h
M1nYn75LZKU8fVG2Flyk9HfjLuJMIIqjuXFDG7Vz0fAsazmkY7C+6oDQ4hOunuwZ
Hczsn8h1k+X/gWM+g1lqiN1Q+Jzv9gFmUusloCZz+QADpqiOeeGPDYbiaBPXk2Ia
iE1Zieb73Bn3kf8cHIRMxmyhcE/MPsMz5IxZGqOtBmiS8zZfO4BHfa7orJzaCei1
bLkpHoP58jN9hzQ621Q/xlXSX7OI9xx+teEpLiLVZo4RKNBU45wXUFuUJJgeSpJ6
l1fnTsgFXolgML4+gQVoJpfIQKiKDwiSneA3pIjHFVfxK7MuLHzvGeGZLU9iwICk
9EIg1Dthlqddc5SqE6+wvL+2E45bDnJhVNvDVVZ5535t9FSWutIIjV0lQ847TiWi
yQ/a6Emyg3xTd+dgnQP/6ijuUKXa2mNUl3kEbz2PnHE7BrAZh+z8aLfOct7oVmnU
WmsxwK1YWjIVgbFA01Qeqp17yLCeNwk5b0MYzQvqu+1EhfJaK7pSDF1rkeqosn04
ArvsnLE0Jd6vzs4IhH4gDZhy/yiSPnKJTjVsTf27rDmwtn3NSkxgRuIvldg8kpvq
DmQ8WWablGNVcRy/NqHm9cYoVDoyRhkAc4a2b5k1JtoBXZGwUc6o9ELVSrlnmWaW
N7+V6SJ/L5jEsquHOMxkMDF66mxojqKlP2k8uVN9wC5weduAK0VXz4w8l14dhx7z
qpffHmj+Dv1otxmWtOuWpCU3eTy9P2E3aJE8jzH34Zcmc8Y5yeDFJAQbHMYv9JCH
Wd0qN38Ldunu/yyEl/cCOWssDzhjgGrrYYinLk5Q2puy1sbhwe7qwmcYm31J1Nxf
oTL+DaJQCXoXIZZbqC/Z3T7DO7kFugf6oINQez0ebH8qQtUCb1/lbaYhHWrS3H30
WmUNDDDnoCI7UX9ZEIbqB5WSqImCyblArNl13aaoIp5RoJQ58L4CAhkcRpgxa5oL
uvedkW9hTTf2sOKtYTBZ0NGPRVRLCVmox242+LsujUAbeuJNc5Ecrb5+b4MrkyUX
4AFAwF7Mt9T34VKYkauM5AicOPM/NvdyIsQfR1DPO+ClmtqC5y/lJ+4vEfGhN0O3
kyVc97QaVPQOFnN/dQhesCM5mkyuOO+TptGIHfpH7896QKK4GMBwycou4SmBED1x
nEgr216q9aNDjcbBEMtmCJzc8L5Ujx2MmE+1Rc0ww+0WxSfrjdk/Sa/BlFdK/AbV
80L429ak9IufelWrVj7PCj3qX5GAJOKQrbryajc2nYfyiOWC9JmUR3/12vqKBUH+
DOljzX7FP9fjLGZ4Czgp5HjGeIFCPxuBzFP9Td1e29g2qMB9R871kY5WRmES2N6R
Tr2Q7wjStBzroCqFQpnARBRYNMd2YmN3q3BJTmV3Bkmuyk45aCZc+ulgW+ZpiGFO
lBidAyzkbktZCnZ8VQYJGvIXfwToUJJGxC3bOr+MDqqjAq8gF44bOgCwTm5Jr2P7
fLKTVysnyarv6f+uIew/djUjLztOqYhY6asZBXKrl0PU6mndoPDAxT6TJ0E7Vo8m
fok2hkoiYjKJudqHcpX7KO5SQqNL2d885WUEh8reKcCeCYcIYApqqCOyEfPkbbVo
c7lWGVtbkw6zWAdjhWD5nK+adyEmwLw1eKOkxCNeu5g9ZU3AqdAvOeOQ28AJHDD3
VEx3SBkoaU8pRbsXwsegJwv/+KukWWX8qZR3cgeEGIOph6y4jJkWNpIcpx3ihJyG
J82HM2aPQERLBht9qIFuf/WgMw1Gp6eKPFb3hNiebSM/7WKURD3Ch3ha4VMLfhDM
o4CwuZ2RG5LERmbtlzHICKw1xDVAiLuEzl7TPORUpEmjM2AVtETGF6GnncRcok9c
TMsdpN+ESYjuSsY3kdu8q/OAbqTaqXe4Z+8wKTckxatf374Waf+3LA8Nc2LP9eQ4
3+NrhCTUuVk9DJs/f6DSJ8wqZK8h3uGgNMqDNIBJE9ymNBONenP/7KnEm84v9+R5
xncwrGYXvW9SG1fY4NSEV+0aR+2Fo5oBd0RThA54Pg0W7TcuEnjrSIL3+2pf0Hr+
eX9/uMlMQXH3cQYet7lV7zKWNQ7cJYgiVUgutqAkxxKte+F/1dYPRfQhMzwPhuER
ctiRCnTF2yMV4e3GTDwtPC5spsrOk3rqxIuzjx9ft0FBYgX6WKuORMEX1VmEpYbe
AoK+FrW/kFCvKxqUT36DOKHKNYtC+cJmv/BF31Cl81KUFxSqy075PYyf3KdQlj2Q
FZoIbYYgNIQp3GRfL1ArZMRGLb0BTsJGL9EvhJMaohfkg53Ajh/wVlUx8CyIF9NW
Pp4P8vhQou/Ibb7qmALFOXa2cspBCyaNBBidjxS8L6LqOp9wbdVxVeytIjzRMEBu
V2wF3ArlDMne1fixT8adA0ggqM3yyA0rfWTAfmoB8Pgl7ikG/KrcDBAt+fQga738
IaCsQR0+5PTu5NRrSRhL/zMTYAUylQlkiDEs9h2SzYWY5eucj63fYS0J6R3Ua5Fx
TRs/lzFKur/Hfq2GlUSwvd7WpKTLHBMp/YpaSk8M2m01RnNKeq6qN1HjD00/AjwI
eWA8F0P876SvRJ4JP1k1glZdxHrsJCD2S2gfaEGIugMAxAGvK5aS4HHPwfGOQDmY
jKg9wwc1R54txPM0k57GPOkv9jrmwkkpo+XHW8HLcgg7MNxhsEP+HmitxXn+d4PP
IJBNf91ZebPIWPX6HX+9Wr5BRHJ3fcnsoWrYs5veq32V1ZOzakM9Mz2rIpNXT3oN
ejgczgGpVLX49qiJ/jbLeUuCOk4NXljraw7fbuphPLkMslm43fhJ9kFBLsdclr6T
lyqO1uQz3OG39nmTl5xJCtX6pCC+0KB/RCHunEugAPIjLRG/DtWRtTzIatHUNtN/
rCenqhl5UKMXdv1V4/LLxxtKoMVptFnXEeHrj5731MPGA8YFrz26emBt7DYsucwY
QisobapeL+S53Y2s1SFBG0Un40+XLBHmvbetH7oQEEBI9jzhJ3jSfEIqwYF+5d5M
5BuOOwA9q0JxwPjsiC9in0BVg2mxcxTgugeOualBCpjpHvigL99kdwhI3xVv83m0
K6+r4eriHpQnuWBbQ1KvXuxcqQBghHAFWYsCbINLKDPXEYu4QBDipLmPiQX6o/Ij
LehulXYsj/UNWOdcM2QR285G6W5YmApYJK04lXrjogoHwyn5mN9DIZawCa+HtLMD
m0j1SQnXCqZKznf2QuoH89zNYZkkC4Bvo7zRdmxPM8GB30CE59QQ0++gFfYuiNml
3NW2JtmP1IjXf7lhKwrbZjPLaTFi5oCdeqNFfojYtSaztfTPEFdAMfpYlJcVc+VA
a89zPUZ8YihNmq0dbTPk93jBpaZFwtko2aitU3EayC7MxLAfWHWwc/cU/fV4XhEf
+DtCLxWSYOzSHyN3qldfKDIBUAEelBq+0S2uEbbCHzVU/L9vo/9ITHUzD27rY7fi
Tk9e/WeX4y/qYzHJoM0vfTwHUwo+rjy3qctAjUPkWVIXAyFbQP27UudxTZD0sKmJ
kmZdeaFycVyMvIDxTejjHxUvG5ihhSUF9UZxcdf+9OM9IF3WFnXvsBgZIy9Jm/OS
tZm7PNj+MvCSwvU1QKIyHv2twbIF0b5USN5QHKx/5UCPhkQq5cT6ypznRwFXvSQF
EJq2qYweSsIz1SSmEtBLVj8Hzi69jnS7DgPSmhDnj6AUarwoT9m8H9BKpb4YqH0M
iIvYckwBg+gGzCUOMXaGc78gZXcufoA4w896yFFOIddJfRrfrAfJncf8GcnENs2z
nI3Q1v2RtfWI+2FqNv0Qc0hmuOyNKpsVn0f33GvhdVC1x/32NokquPGqf7lBMBEN
7jaMnqRkv1pJFcrCVvLAfpr58hOiZsa0a/X6JhmIKQgCwcGsZ3rGHXKow9dYr8S5
sce+Br9AuFqW56cTFWqLuTlzNpFmnMnuqlAnKs0b3trpTQdaX13dWihL+0fLLrOA
nm0mBkwnxyFmt8qsgtgwa4djTGqrjuF6bkBxf0AxuBdsjs1N3k0Id7vIFBWHpP46
Y+AzDeALqNrfMpKzkmjlCEPqcvnItBCzrui0i+dw2ViTXHPG/qgaTGMI5HIpNHBz
DCuazK1CHrYTYASEtqMUqnD/dzrL1bhyAB+wGsLFmxx2zcppECs9lA8rMiB2FEa7
azrv+qGawH/VFaK30kThSD0SOgywWjLagB7O/C2B8OFjVhJzhfwWf/SwxgmV/FdY
tEVimyPFzfa7ImynW0YbVA4iBrICppbamHgohIJCwOrHrbjluXhA1vJIbm7NeuQE
xBHa8k8E2yV3mf9oxvCmay+sMk2DyPB4fKXvhXRYwV6s1zsi0RGP6q7WITFmmwIj
aRT1dfJuQjiz/982F1fG3OaOrEhGd10GzYaff7SvZvylJSjbN+Mkn9sFWNYJbFaC
83o1cA5aqCZLm1M5akFPREwvIOz29qppdORshCBHqhk345w2csBRYfzeG0imLqHf
i7G8AH4aCpi/0oxty0fkEJyDQ/LYfL5kzeUSAupjZ0uPVGPWXfMkgB4liUqgUwnE
i5yW5qqZihnxpeYsdoPiozLa0tAZoo6VNW5CqUwxWHsDboIqnUfq62TT9Qq1RP8H
Jts68WgCueATMTnXCq7/33iN+x/5R9g42qmrs8pk+WyWxaRFCJdAI96OV2ya8Wt5
qVFKaZ1WWb3OZCunIGy7ZN0JB8kLakNYyCGKjrwHPk460H3CRwH8a8VRsSYE2iaZ
GI6EUuRb0VL1L7dTh3MAqKdDpjgJrXIOywFPgYFwsmQKv/sBhY0Bg7B/GVA+EWWw
nxDBjGd2IvuaWLrpUTSIRlNzhcQOdI6i1mtWjkXLttMmOsvbP3wtMDuPr8PgMQjH
eYAXCRtE1y5gR5VFZx7rYIKljt7x76Yvs0BTJWODWVr+7g9HI0ZP5vTTWXgk6bR3
3Ec6XXRCn5VE91yixQlJQ0hJqrmqJ+kbP5sQXInONiRk3WQ+64vC7TalCdCUg2m+
Ureyb1ynK9thXRpxqhUGYJOKGZut0yqpGl6LVvotHG+XOwvsaoJUu/hKI0sj3hQY
RyIIt1xgulfMPRNlb7MxzEFo7FikvgSNhDZGx8h+BIGtd8zB0ZDPv518MG+LbCUh
rfhe5dfKIBjtFwI7icaKMpYW+CVJ2qaxh7iJ0eJVNhMMoDYL0JKqXRuvhytVxL17
DH1pqUuM4zRgoE5k7pQuaEbe74dt6xd72dv4mzU3et/qGkjtTseM3nSzx+YT+WpS
pVV02VpacG9oVmbfH+oeZ0dXTV5inUVcawRPx8CF2BvVCtU0KJiTjtVTqPRUqdsS
/v3RJhkIg3Mizj99gCONJ2C1xbRTqLNAONbNoscQexVjwKBcFXwfBv5u+aR06R5j
as+7LIs2N4Xeccv1StJlT7i+Qu4JcunVxk2moRAScPEeIsNFVhcBUg//DgMM9SPN
WPX8NQ1Gyg5nlvGvmCBa0qGlyfVui7uKwXWRrpveMmEwlCqdKG+t6F33SlmpLLPO
40qIkd5oHA3Me7R8+s4XQtPlItUoUda6wmEsuIARrh0y5VkIih9uY7mptMfrcDXE
HHGk70c/kDhtSCgC8OfytOCmDp/cvqophXgvaDyZEj4hIJQqLTtqvfFhVZsUS5PQ
doLH729ED7zzuM5czWk1fQVFiyxr3gYZMHiswoXtgospmuCSR2zfwZyhgl52h+6b
JTa3vO5yBt/sQiWjxUxgSH7rNB1nwrRChccz8Dors/LSlRjTWYT4GJKaUAmhA2HM
5AOOh+B02CQyvOhiPoVfHc0nv1DX0iV/+ZHJA0AbZcGcmp7L8e+DDPfprlA/Hk83
POFkuywz/RrwIYD+UVpnkkytH8rW9nLx/znSKeqYsCoSIuNK0ZAA9jawQ6z3oRxS
reG705dDTSepqOLRUxDs76R1J6Q1cUFPH8kHefdpvtgsQrpyyAjbo6hd2YujZPw+
9Q2fxp5MKoaEzMd1jb3XzWtcM5Wfmi59IqZigJTXwlQxt0HhB4ilMKnPjq8XHLu9
IsA6Wf5ZI/UWhw6qdlTmQDc/cieqSp4toOofg+Kc/6S/+GCj4rWhiUViUo81ngI8
1acV+qdEzYT3qERfoWUR1MA/SoJP1LaiUI++ETAg+HxPzAJHu99cCNDodlzC9wYS
kjpMWLDeFex1Bc6jB76UsacspkMQz8BA5YVYdbRbSIU3Vb2/EfDplDl1g9tecGyb
YhWEltj/eUedaT+cu9D8GabARAV/c3MNr/O1s7L7Zfdlh8wS4zfltWfHWFSOUsFB
HdR/FxVJKwGrv+0tRF5yEB4ZCMqdX9qPq+8kgv+aTtB3cu4rzeRI3gQfKwdI1Swj
BJfjD1l2X2SblL97d2Q5E54Ipqa+pzRYatLcvu2OAxyttxBcAWlBPJNuni3I66qt
dkCkdtxMIAVkxB7xgfze83lRcAcRXFi7OOLa0uADWjSCbgv5tWV6dj2dHPQJuEaw
2BdnxFnP8XaF5c/5eoKDJRowgmgow4MtK8IM46ojVxjuKyY8d+nRaQtd4XAHvH/G
3WcoKJ/Bx8WEDq5S90QcQwgENwKweNQ3KwZkP0gXzPoRaARn3lFTw6aN/hNxQ+zK
OAlMv4wzUm6BuWWwWAdHU6Cdp8btwvzhYmHCb6YVEXckNJE8dW/8YQbbZaFWj3Nk
vazFP3U2+o1T4zMRLwS0xJLnhRQEDlagywfXwQN053HizAWKBMVZOxqTn/BOC5+k
JQ1wvXJagfUMXjJo59/xu+IkO2eDd+fYWQnQ/Ume9NmUmmsLS6EShj/2tlT8kNJz
Puy7tr+51DqIgavGSb1HKky45J2crz5dTElA7A1MgeLjSrUA0PXjRUdM7R78HSSb
XSwwUHSLY5aZuvEADj4xWZHtmpfi8o8uEA4s11A32hcObKt6dVJrYC5wTLqcgsiE
pvkY1L+LMiXKmKMtQ1Vj7neOuUOrTi5fSU00W/CiUeW2KE5lPP9PPhFGERUQSS9G
D19HY6Ul3FzqalVHjasIEoOptFJ/EFgf8m7gUXaCmGcv9nyrgSD+crCShrg1xGXe
sDrGgl5HSEXOOlaNEjbwe1uY/qL4vqbZH7WHFlEETcnW2Fpv91GALmwRUrXHKEuZ
1P5Rq2lRHICVDv57pfDTYIckUhpThX6ySmtF4LadSrNj2ZAmMPtMLcJZfzlkg+1T
rrVYOU4pOE4/D6hJO+kXgAn06MiA2N4hD9t/9WKIvV7EJVghAPpOo1D6HtFJQeof
G8L2uuTVQTcJsnWE+HGRe/ndcp2XfnY9pfFXx/SeEAO1+JmxPeT1dEOX251TQG3i
FSticBR8c3imeYQ92XtuMtpCLHm2HuSpUreD9eHnoKUYuHIIMDBAfUf8GMI2SmM1
QxTYBxYisef5CVDyR7ISMFhSI65phsS5r471R1ZgFhkWPmd5J8o7CiR7FciPQPuk
ibt3HpwKU3KHBmHUKuZQdK4URWehmlEc6IhdUDALm/c8wH344GkYrUIFZ6c4K36V
tq9D8AhJbQnV6CxcaXOEwVErmCazBx+L1V4heBn62MF4UgfG52pj12zYxEH4FqvG
cZPGCgtA5EyjgmTFCyMrCy0nRQaWZyPzoV59rbKXtW+4ce7SlNRQspMtjPTMHjDg
OmQvmUcBvsqpsTN3xMGYhhj+7cjuTM20d8ec7RyZAzr/gLAK1ALkQxdkEvZlIRci
hVAdbtvqzEMqwJ1DzpEbhqQh9/vqVjeb0feSKoDIMKY+tgieL3rYZpqCNiOMK4i2
wObHNeQOiyYrVmeoYZWn8Q5og45jd+fnibZUP2gc4YJvwP60bs+ey5VoL/Nu4h/g
rAQorBlcz1WdCN3gd7nTKfIuJPTPqjStoPQNRn4rrsOOFIe7d39maYQljw9+pdjV
cmXFRN9bfVnARAEr/09N0H3vDIX1RbLVyBYI1MFGfM2zWOfh3ZiTOMNxQltU1/pY
1K7JiY4tGyOR7CDXUtrCWVGdFR2c0/T0ORVWTc80W/HY62Xpxr4aNVZpF7ZsHP/m
ug8qhypa/5yEMi/2w5+rbEYNqc9pmLQVP+VexTvZL8/a9KUM5245ax/Fr0e14BGc
7zl+FvNDS48tlCw0hdIUFsy0ytw7OvpG6p2wJYuIXtpuUYGeAI+0+UQchBO/Shg6
Y+HzbRLe0Chin9L5sV9oO0jGmwokH67FCRBPI2GV/uDfEN7tPy0IAckQa3wgrP+G
C1KhJe12m24kL3nLXHA3vNxmC1XtQvbl9VEIiqQLrr9d2kcaIRPoDbj5pXosYpez
cSFRDBWiiUf1JV6HPu3u0wXIrccuLm4hgZ5zYTZtPA/aive2ajDEPl/0zI0tVJ3B
JeHFAUTFlgRLaTbvToWd+lo2YECqMyohVvu9cnbiHybuP013yLAJr0fa5I+QAITH
bUujaSuJnGoszyrMH/CqSR0Qnx2bylE6kixKjRE5HH6bFbZgx6L30MFAscMeq9Sl
KhLS0pNrWS7NQSiB0HpUAmIBbhCrgPRZjH79vhUMBdHKyRi82Mw44aKFoOR+d93U
JWBOKyXLgeiSzfNpvR0wGV+ielsmNoCQcfykblXxFJg6mqCEsIQnNnlvtFmMk2uG
vbr7e56EZNY+acWnqp49FKBQBkuB461qp/M+EZXy2m5SsIMqJpOicjoitA4zXUbZ
XKzP9MCeT0Tfe6qIZ79WliSbO7Jj0fR6He8o4XErBrrDUZlEHlYZH1OCI+DqEcKl
PyEreuxpdGHy5BC9a3nzuijfpgISvab4MyWslGFaiZTykGmROiUwMFpIj0oYo0+M
1VgoUGJsDBlsgcd2Wxqajt5Rke/3xwCQUwFFzSqtyAELNwRM3elCNBt9QruOjMXZ
fkXVXcGjOD/34qicU5IA6RhoKBy2WuSXxdW7wcqWB7JHn1fLCk0uGv+vRXUeVKeO
O+J7qb3YRbhwa4P2G1DuVNmPuGLPfZ7un17c9hDah/XmWsbotxGoyLLdcgDxrrwp
oF6XZ9l2wUxw7cQRawof7hdiyi02Wjjie3lN9Ol/riTnb1VIf3BgWq4O+ShvWHgm
S5ZAQBJk9ghtb/m4voQvUI51zJp5onUJhKgkIfiOQBQGHkCw/oalgXHuL5soVjOU
DabiZqbH4U/wmvOzIAw0aBleIZYqtmXQ8YqCIhTdkp5sm1gbpRnWXLojMmct9Y/0
BI4a2FE5noBgYEG96V12YDDwEAl/bi6z7toua87vOMelKxaJNUKnwQjP1Hstiiuo
xXu4sC/778etXy0rkFE/3BIZwGT1LPFpiOe7r1dCAOh/36sOfcPSt8RHxMLHhEHX
VlCvYNNXrmGc2TI5Lmrf7LZLwTsREgSk8EKkly2fYSmzk76oqP+1G1I7sJArtq8y
K84FoRmePp/8DFIfeVfhl+sw7ePJ0A66M1vBQy24xtw4d9rFQ9oFSJMhs0TqufhF
Tm8SNL8eHcwy+c7GQAaAGwt2uaUD8RNsZ3Z7ig8it/Yn7Dski48G1aS0e+7zO953
zzS0lTTyBCB7NU8Shzd04so1/+IfpkISLRwV7y84U7fXh5ODZfrpO0YXyyFGWt+w
Zepn8GYC2uw+iIOYcoxXCRGf0L9c3ZSwYfQ4cSjJAbI/GtTsv1Qnzim1qgYecodM
KAjrZw6/Tg3GFs0bTiFQhnpnt7qNsRmS5BM6FR3xDUkK5CYf0eynnGt1zfR8yxqK
jJ2ZhNiBGg293MkNwleJb/uhf4O4iNckRwHXIlEfaAmfhp2f2zNWQooM0l0UUq2c
9EQOUODXdBsgNnXKQPPet+8N4QDbJsuvMWJEBIbNtQPSX4iz0S6BvTVdk5W+MHum
pBkc0LtECo3UnT/SWIgHAB6tnCF7hNiWcdQCL3Lv7nOae2rA2OPb8F/whlCsuqOe
crbn6poL/mRqXRQHU3V681SzJyZWPWRHRRE5YKVJ0i/4GSx5JRpnau7QuljFX9I+
//EsUfH5+vd0J+lWEW3OIz1KLl8wy3JHJOKBTthJc3Ks1Yg8hDSDEQaS7q6nIFDA
2HpctFEdMqCsKNXrJeQztkBiR7YGn/YCI7xz/qdtN3lV24iJtExmc0Adv9Rn07Uv
sk++tIwFSdftEuhSu0GQxfZe3OZ/L7fZh0Y7HOo7/p9W4yl0J5DuvVVtqFXDxVfm
Olz5avynHdMJHKJ60pmgOuRSSfXDCvcu45tNefAdyfi2xsSsinb9E5OV3Q+pjnl7
rdddrYGVNYmUwe1ifmOorIYegqUdlkwbTDnfM4jbBm67CtSnth0U4YvEcWqCKufs
SN6I4m/CWTxKTiFLjVOvrQDJniF6QMIUzoul1neW3eu5KPq3GK9c83WREJ79xcDq
QV0tEe8aRE3YY7keq8WFvKBMUdbdRLYrpXVHuKd8TOJB9miuO1wu2Me93ISTPBHr
iqmR9iZ2SzSO1nXEX2lAEd3lNRwFQIq5fkTv3BsVffFOKRAAYYL/rEo2WbMI9owm
QSPSYMUzjLVr6wBp1FhBKhRyU7OOHvYZdIJIz8axpaxRdG7bIZ4o3mExV9iv3wba
gjpBwcb8f2FZeHn0pgDd1gZOqLnJZB3W+3NWaLx02Z7I97aXotKsSTMIVZzxWk9B
r+NAndv+3i839CMR/HDuxPmp+jjdEbzYCyatjLxPQu5vUc9mfdYi/yaq4sgbfXxB
lL6KTit7bAsMZbEbpAuWANHItK/8sVBYjdTVEquOXLG0VawoYorYGOyHQXenpIuX
sQCfbXV9Ksq+BNZgYv8bw2ZdoE9+4fXoa/ZycU6Pg6eDjoNVe1VaPJvqnvGGEeGX
2+E7lPFOijXb9XYpeoMQH9TB+22ylXnMsPCRrtgz7Tjr8px2Jzuvp65iOgPol/4V
QKveBMjdlU+yKesY4rdGP3IfoSKaj9GdtwvH/gAyxCHUP4VBtRo2PZGxtJtomvWT
/+Y8trDyUJz+ee2Ol3r1bR+pFlg9EqFj41703xt+bvtmX83NV46g2TJEeGS6BCjx
jl2d79W9Bq/si2BOaoxtX/MXYC4jIVZWl6ypaRwn+YHDKhw2sXdPA9G2Oeb48CbF
3t5unSRegod7ooimnFPUvKa5PJrU/of68hz65dlYX6pkTa+h54ri3dWq4Fy6t4T1
SZ02VQazMFwORI4In9skHiHngnbw55y7BEgCXN3vUWK8wjJRHYyS2VNeOCmyIeSq
MNQ0TKQ6NzXmwjU9COW4XeR6pFF1nLLnypQarqFk2qGwKeX2Zww6XK/F6LKX18FW
2/uI3KlaAJacYAD6hx+qymIqkZAR78ntrXkadlWAg9qBeFskeQ7VcRZLWDlwnkUf
B8A5yA+7xSVeCvsaaUtdakSM8X9Ue6AKLFiwvEvozLKRdHXSJwCyrhqLRK3appXn
VkHvvxE0Rmk4My19MuStEuGJfO0CydLmWFAkXo/BZxByxkeyx8UXztEEswF3/cQT
4wbaooHnhe2tU22tCBP9KiCQEvEkf1XVifEC4EcQ/twwpsvdLv9t+c155Hveb4es
g80RUWEy2kyp2O6v9Wlrr+/z54XvhUfY5XcDhWC3iv9G++QTl+fUhKhdbMe3NDpv
zLetR+DZKpY6aai9ahlb18zWP4grLMqJN3i8sOTR5Q6OEd94DV8EtKT0vvr+Q6yc
1bed46l4xuuBsunKLX4Xyor3LqmhB0STW3KZOQQxvHH7Ix741QVcR6nd8HbcUc2C
EyVBzulxx5B7NcqwqSLmSLWeELtRdHvPv0FpeG6ioFDkqjRQRauOgEhaMCraltlZ
ri/mKxRLUg/NubUXpIakifMK8E0HF+1GbvehBOSyUnGjtIZtj8fIv+CtuiWM0HT8
KWCgt/HD1om1+z82eZVN6/fY1F63rbsnBXg/w/zEKn5Y8kfAkNAexRm8/8JvoWOY
bCxPnV+fUkCvBNK+erlMYpk2nj7P7DEryYQ8ftgnS3VrLw14YgVUmni4VJ39gryt
TgD38oVlPnnhxnrObLzFvq5EjCk3tQFBkBVCA/CqaoimoRMyIYiyUXy2l19MOWsA
zd5v95u4XPHjtSNMJ9VgI8ZB883rb+i5GPRwqLzzJUoF0tB/5WaNKWaKZRucL5Gc
6kLcrDPG+KJ8pefqJ8jzIDQk9ZptdcqpCcxUJENNFx48o4J8j1+bK5SWJsQKhSKj
lR+qEK7O9HidSumdYBCeo0/Ow3qpko+xFpJSxF5MXW0ggxVL7jTA7CfKUrfpGrSk
RosvhY+JAgXoUUE6ZwA67jaZNhCoP7S58S3Gu3xIQlo8IazCRgz2vp+muDmaFvZf
/EVcR9qo+9iz75HEarVfej6Ka9kjE78eljvM7yOkveZeSbyqfshv8CA0y/o1m546
Aij34/HoNSFgPKjOJHPP95CZt5rjDnC9VzT8nroCWqIeIJfLvlyBUldljV2MTrfX
y2cGvrYw1rNTzzyQTfS+1Y9jCpUMh0GGZKlj9NstTQ+cOzmfEF/Z1JIaDa7VHPSc
CgZP9ODVBidJGQ2SEyUnPDyq/B56/03flPqbtHF8dRuzLHr5WSsGePMHVco/yI22
A0ZYpR+UAdzYVWgxbyCISTBE5tCmOaZDy8WyQ6Wi3lkK6Ez5TsfPlHfXgFINkESk
zJxpOxETF2ENE//Fq+59zWTJ09fEVNgSEaTglQRcGeRPswqztG7JlPsrtFCvO62D
RYbIjIW6wL204ZnOouQsGdG0TdXZw+0R/LvyXxM8xc+nKDsUat7h/ioZvPHP2Hnp
BrMGW5GIOxKLIveCcr108fGY5jjbEq4462jfMnM2d0MNT+4iGyRyIsK96l4R4xfk
p3mOX7KCDFP4NfHjRwZylQ1zpWPk4JD47/hsmucIO/inJfYVTvCyoDT7IimbAnx9
4FAbkD7f6ToFd8IQe1P5svwGplDTqLiz1gR7QQtpDDGf1j494myG2InAy4GHnhz1
/zbhLeEIbWiqs9uXBkXHCvv9XpkdFqI8469CZEUUUBfxNL3puBMHnSCRlavKSYYg
k47Dl4L/Z5gkxDWAtUayM04npi43Gx9ttW7rgbxy1OkC1xAkHpHTEw43uuAXSagI
4r5jWK+QapsKJ77kQ+uHD2DdOPnZly90yovJqxhrOST58BcDC5ww4JCxU7uQdm3E
MBQAEKAh3aFALxQeQdE48ytmgjXnZ78cn9tez/pSU7/dFsyWso3g/0j7b1E/HcEz
F0XYO9SCtIo8SPDya4gMMDWj7x1iElffSoicOrXZGTxt3DMOQEednIJKJj2UohtX
9uoLJ/iUbEe7MrVzEdRa/sR0reKKEp8ivOkgeu/0FZCV8dtOWAOebxHPeAcEeLxc
zkublfVHIyVBPnhy2+myTFu4PopT4ValspHrTArGpU9ZflbL4Am0cI9qJEjWGexS
X4fEH5lM7fYMT/T4C+dSFpipkL5fU/uuFUmaShuzKPLE2DNhZxtJ8yHyaBaosYq/
uyTnTqKSDXRCww8Ta2222d830PYl07YhqVepjI42hUPi5f9yA7MWhuUqtKDK3UtX
THlkX0zH90RNotmEymrRV+5d6Zf7iKWcp57V2M7wGJrVucgf2HVWeNA03CJta4bR
h0loY/opVjklFUHvm8TX54x+es527ZNoICMOZjAfi/0Slp5+4yCm1Y1twhvYe072
6G2mSrRfT3hMaoRbtFTD3D/7DuQpuMAAxxLjABWuz41sgcN9N6dmTxM2SdDL7KJH
OsPxoIiJIYY/hwh9bmliT87GZiqDlixBDiCLlFsnlDHAqazRC0UHu/pIi1YqX5SB
8d4yhA97Auy8yLpI87d7yJVY9sTqNRjRRUtbIxhZynDYNyQ+f5QOnD5aSomXk+mZ
ZkSaGByiE22ArAvaX70f4RZUqNKFEIyvQ0GoWJWN9Y2vzdETA7ROxqu75xae/MrL
IMrXdthV71wf6zjh+TYyAGEkOdmMmOPyl6xzdSnJ/37KhpwhM9ExWF78ZAGaYg/8
yZzMu34IEwrcPDRbZ5Mr7dyLUdq37ZqDDWXjSc+mmLuzK9ox7FYt+IRT51xWDMz9
CCw4b4TesLgpLIofWrpqNI2X53IXYO+/pgyQcxEailWctLYRFmHTEo/Bfp7ZcBJ+
dqkFJawvF7qHeGgf02+RuUXiBpRsd3WeUvWLha3tKE4rqC8b4wH98rJ1dIq/Zn4t
0bkxn3FvE/HTLgxdH26noos+JHyGKNHs63BDNmWBNwiFyJ1bpO6r5XUhdF0dbW0I
hhTPCcXxrKSmVtCRoAhUxVcSTR8EpywPk1voul3CF9be0NovRvpH420lXpn0RN7k
un330uoBo+yRmKdqWkLTiylSbmtS+FyjGm4EPRXVgdQgfH2NnrER0h1iuMiPKHUO
UGG2sQl6ifmRS24E3vpNy5ZTHESU0WEP3X5lhY/cPF48t6KYmsTmLOQaHqlYqs4F
f8ItWJKCsAFK+1CgkOEqSxRc6f7TqGq0+t3lsy3pLbD+DYIbnhuVTSGIwMw6/U94
sP0ohjhym8jWxHcUM7L9mV68uvr8cRFh7xUO9QQFQicg60W5k9p8xHMhrvbMUi53
xSG1+kd55nKAbmM0X2Ir+Pq1bkiRR36/OMMnvDfNQbb+RxRSmT3YscegDfKcvuFj
WCdxbhdWFVqR9RbBm8IsWAfFYW9RQFJTb9ibUmvLdMwip8kk5URlnf72Q2MaVoAo
bk5x9GC0FD5VVB+dzH/dNsT34TVra1mi6QVu4Tz8WgMQlY7mZToiFbajsLqU0Ay9
yZGz9PAy87du0+R0DRcJWw3/i9UzjGT9uxb1sI+nORfzDQ0m57NNn4epKR0cbIYj
1tfKRT5SHXV5PU0CNWRs3gYrcLpWFrgTRYqGeYHBmavQTdf3smqgVfv5vXp3G9XB
Z9kd6CyqpBhKiZt6uGyLjL+58RpXGbStOg+C6VGDkESSHjTCK9PWn+LWfzP1T2dS
Ra+m6uj4VGnM1I9+irA4FoAnIYTaKF8oVYUfMZtYIVAKnYuw1ABroEwgWUaiPmY9
9GxyszpRp8Eq2s47Q1V7XnpGwzKjYnSBYQrZRLGfkzGabNThCYTBPARndij8+ko4
Jfc75R9sVIoJuvHSTjrf9sQ+afDCuyj2mCLnM53l9TePU8VPPqhbhclfoF2iofIe
wvxpdCfmJWfJNMEeepZqSRa68AxsKaJZbdn4lJ4he2CkiUsnLhCC1I9tMsGhEWzk
1vOdKQij0zwGwIriBgwiXld5HqNTKJrUfuDrCnsJdxIETRlTFFe62KrmFx9olcF8
mIJAbB8L08o8bHlI6OrX6BynsAzFzJICvo2H+flQMI8JH9b9WvaMgfHcvIXLP2eC
rFZ2QBODd9tfRkXZrbI8GYjkSyN1rlSrJy0T4HetmUbJQcopG1bwmmKHE1vSNNLV
TSI0REJCJBQZyXz5g5S0/UR4v5vvvhVwpPyK7Hx9XybzgAyKxDgUsHGGcd+zXbHG
14fZJcTibGpxQnThAzzFWWVShQFFgFi0mw1k8xRfklfCZEJpjqaufOrb8vIUKfZr
LeFtrB5t4yAIh5PynLjf+H00YeuGBkd35P0bTVOnFhiLczN8esf8MWP2KqNhc7/+
+jX3wmiUc6kajNlW4PjHLK+twoN5/HqZeeq7/QkRG+USCj+SQW30fblOjbxCDTlo
15EwC7T0cfCvubNHzNOoYadxTynhUSuZ3XGScFyrJr+hVL/Bdjbggnc1nGvIFChq
nuXdcHHgaYbXKqye2hoT88cXmAmfrSIWSP9/ZnQEHYWvjku6s3xFX8xNMxLHkaTK
Q1FdL7MstD9TP37EiNTmy1TzmBLs3mum7a4E4GR6TtgNBjkDD2lFST5FMpHECG12
uM79lj8acNIMleEOmwEy2bfsIYiXfSXAVSiMFOxpDJlLyRIdgFqnGJD4AArIXDiQ
Ty1QVidDIyZ9VoZPrkH2FdbDVvvqbx8DBDcK6Hw/jwLgPy8Su+i4FbqGnGqgeOri
BsKUuKrwW4B+RS1VNiUyQNotD71zF4lmhEOGSUlRNlyQ7VkJ76QCsY/wUhsIeWZY
488/wF0NXWq2QubHSXxIIEmFeLGFwooCKwTvqtCpVNWrR4Gx9K24Pnwid7OMvAQM
EkJb7D4Dh0+s3lMvELZqdV/4J9GKk99tq9XuusFl4PKr5Sw2KOGKJUikemULQydh
H199s7juhDQ6Kb5tt0O2B6VsFIGqp4phxsgCXVRL6OvKK7rskHGyLi5ezkscdW4W
BoQw8+ZrMU0xo3pk89BMsmHz8EQhcT5Vt1hX8GWaJ7sA5FjWoIGzTa6lhPcMRgg4
1LSTgAzcA6Ye47kGrw44kGSkuOp/z2D67iSJ2Z0BgXFjyEEMochCjhlNLOuN+mE9
poeW+N04KuzzJVsRPGV/NHDh1wvvRFglWW+Prhd9GLJb0idv/MSzyhbXvrgAqQlX
gtCZi9x+EVwTXdbgAyeq7tP4toZ2FEcppaa3zDbFbbLzGNHo8wJ2VUbswFevdb9k
3INP480Wzw21TYmC8fUYE1ail9aoalj/wWVyAzogHMOzzpG/+Kh2DyjjDJZmVbu4
ZUuskp4QlJu05Snl/TE6srl1r8KTySNELm6DSdTc9zspzYdNX6CqtSzOW1mW+/D/
O2oHhr50afpZcAskhUCeLzqs4Ue1zmfam+QkNt3ky1JnpOrFiKitbFF2T7Aw8RUr
L589xI0Oi1FEAwjs0McbccHN52KBUlT+m5e2JuAY826atTw84HPGuv5zTnZwnTMx
2d+iHv24DxwJzuY/F9duFhgtPi82CQC/i8Tt0bUB2BPr3tPVxyGwiXSGvMXSK9mM
5Z8xNKuFYxW2u2fq3jBauB8Vhb3zpu/zNz7401swEOOIqDG/AxzBbbPzGRZINTjw
I+ypmw6WF1x4aj8qYb7vvHp0zBrY9ZjC5kJGT8SEqdmvPTZ/2J/yIZoebShqiDGe
YgoPqeMzkQU2ejAYpwxPAZB/qJap+GH2MebupodbALx9LvQsvuApIIt1onxxWBqj
alWjLYsWpCJS04cpivLrnOOJga2AvUOoshaUVoycKRvNyOh+62TyWBHZ5OJ1iC/q
1QMCMdux6JlYhs5A9ASFvwD33lVLNt9Rz4tdTninB4TaDnSYzCRnfIoOKuzXDEiD
lCgMY35FLg7sdEjqZgdKCI6u739rll7oSics1MKEbua1DoKHt9QAcuKBJPSiRh+m
tWidc9T4l4z88YULAz05008/Wg9LEs6WDYq8Vk0J2x8im7YaCUEbeyJ/Ox2tvLGG
G5rzmU0pBMWMs9PMSiZMlxkUoHgz3exNnB/bdFKxMBYxCaDITI5RCAfwC9LLtgsK
Hcl/DFMEbeq/CjELB6NCpviLYGrok8/lMRWISPccvYm9e2awGY6yJvj8K/k0f9N6
LlURAhPyCY/w1hsStOgw8ciM4iEfsiEzrtjCsfl32EJ0eD6kAzSX7sFIzxOLfdj8
3asKiNye+DbE0eSLB5rmhe1vGUQlvZvpF9UD2b/9ILIlh4zZ+Oy5gaNOymMi8h4z
bKSbapWzA3HBablwTw7jbzF5e8iCEm5AiQNrNC3UMvLKFohMI0Vb3oCPA9FIko6x
OZ2VVYWZq8DXlFBmdSL65ZmBz903i95MDRu349vun834S3Xa2rDeDU9CE+4vN498
T6XlG93mVEcejE8Wji3hJP9A2nAHBraodKRohA6rFS2ITcBToqIb139OHE+RD0OB
/nSfP8fpLPXp/d0u0YEYQRfwpMx6eVuO+JbzgKBUSiHbV6TJUz7dQQhngm5iq8um
yMZQkMIKScL2IPtDcDbuTkmUorz1yX3cDNfExqaL9Tu3iOjgt2sECspFkK+FELUJ
Zup96FUo2HCcvrgWOuPqaR9Wg/6719Wqw88ZVOk7JLLEoMDFiEIv6KYCrDYl5JEh
TODysZejHeyP4XOTSF0yO/UA5wjhCVTqC7+cKJe3qi7/vEKkMyFPjjBMGJkWdjHh
gVMrioc5e/xBZUF52AJWqktDg+UoaAFTioFroUusI12Wm8zQ80f5efKzNDjJ8mxu
XZtLhpJkT3jmCzsYkfqkRPFhxSRrvOF+S5ABuJOkLW9ZraXYI/Ig4fu4EPi4iv0/
JhI+9VhlpKXzkQkoBUDlYPur0PY+r+ShbOGsGXxVq3sjcpnAn7Qdb9g1ax3ji791
L8nYHJ3Kf2Xcvd0LhJNm47dObfvPSR3AiS2U/iJqm09azS/7snl0Vf2acekmhyaI
sFF8rc7XDNt6KoS017QlrSIlbu9QxQdmcEHK0bj+6Jdqj9KdwCh6RuSgQ4Uy9nLq
xVgzDhEBBkewwQi34sdk5Od5m+pI64PdXJwYTLUkA2AzacwH41tazcBvIxwBcBD9
Hqhpbx4gmokT+IXndPb/+YDKfCaQMbIquH2YVRQJWr7NT+0Tl0joPyIcAl9JeDHF
iLjOUh2zft4OCC9GG0rGf4pIQt77qY8rTPkFA/vP/5mlhI2lNQFd8mm5321izPbh
VD7PZOgWTbiRViRckxozw4W4WkiqF3v1xVNCGzWfaMARqSQl0Cf2RJEv/eBpX3Pm
9zf3ZUEkCzQ5FQh7CMKOSq1C5QAO75sYjv5rV+5sDdww05k6pIKZIYnVzpfRnprJ
GjQ3tOuGCfdomNmEMoho/1hEahNYv+8nk3P8AHkCKJ48XrNeIC0fvfIRz82tQJj2
AQK4scU+Ah3P2Ito0h1EdCqHa/mhmwge+VSt5zUebQE4KCgL9TW1gAzwngCzMtM/
EbGcH5JizTIh4atzEAZlrHNVX4XrMzAbLaT9DF1oT9SLAg+MBIPd0xTyAh3/Fvdb
GBzpEgghGY5UTTaqvvagFsjgMrHDse4cdbQfy6BMuHW02nT3vC2rnxSqge56k8Xz
iZB1QYlWYopLPjet75sL4e3/JZmPz5XgF2ujgYs74IQaQStwiYcqpMue+OTrmF+V
cxtds5QAEs7KLb2UE2gzuubDm61WG96AODU98Xx8kmCnYCZPMAEZeymUJ/VRPNi+
UZHEHdWCCR9sv4gLaIYkm8injHdn5eq4Bc2QaOO/eV4cNmHFnHW8xchHs5AZF4Eh
muSvfE9M43H8vZ7MPpLab+ERtRZRUlNDI/3pyw8UIABDzBWK/qp79upj9U2oKx57
Ht9KEwEZPH2tb9judvE2uCbLNlSKGSm2poxDKiMczAzWhZsTuRefJfnDjvheAFb8
sC8sUcB4UTvx2Ms0onFFXDVuxZasQjxPsbCCB1sgGfpteIUBv/RlXeF+fi05v+a4
PpukLmr0nZ70eOxfV1L25uAk9eTliQA+NaArbthWYSpltE6HbhIT9qtYx5B/kTHG
DrzSt+W7X+xMVM5ZAWfAvQN58xrbKxRF17dKSOgGQT/+iHvX47wiiOTq8l8C7rm1
9XB8fUryZT2E+WGwH6x9dW8ALHa2YIwlUT0uLBBVXg2RyOrZxwZNxUMtJFNH0eGq
09GgImjTx4sg22P6tEMmVlVRPZR/Ft6hZnDI9s0MrgVM/rN2XA8qQTUKjuX1BErv
Oslib2gj4yzczXNMZl52xhkCEycUoJrURkl7c/mrNNS+1RMlDaBI9NI6PDkudUyB
/JU8zANyBYspX5GPjKVpL6xTSdd9ohGlw/zq8KmE0tPOh/GD4Tq8QjoxBVAAjYRE
mX99R+ib26zoA0IryvldEKcEeKnoVSluiM+jJgr/EOY7EfGsJokDq3nd/2tz3mPn
IF5T2s0X7Wa5Gekuw2BF0OXYG7hIB0evVXzcKxk0hQd69EZrklCorjEUg3OqzF/C
x1qjOjOQ34TU/VHAGR25Vf4x+0SxzIT1kbLXSrsGJTitDNBpasqjCTpBSH3r6F4S
tON8tV31GmhPW8T+IQ5CYJvK7qYdYkSTYXvmieaKct8dVY5FwNltcHffzBofj4YY
M9l+UsB7nspPrxAdMTtEFQ+3kkyLGCVKexWRimbSrkUUtkVyy4qFb5ZFNFOrHMmb
1OTjqGEmdohr3MNqg71Hwje84tZJJWG1qJUbapurYZMVrHPfKgQp6o4lAr5vRbJ5
Z/zK+CABxDiJfypG80KEjRBwFE5yueQ1oiAbw3cjE7+rCPzlncO2DGKRaKkFnpQU
Tt0uz7lsyIWeV23ahmNNBOrLcIHl1Jq5dGtsUvekTLjNF7D0uQD+fXiKlFSRTnV1
4iHLkNwSZQbTjhiwKoN7MkpDweTM7WtahHq8nr2E/3N7dHkJb93Tydwb7Swyo4iX
vO++VOce0D694mqRGQzKXpjggDomje2NEy3vHtepBhWgj+xqMxxmNeJJoOQ7jhf2
QW00/+juPPZGW/7WJcYpqq1XmIkbhR4DWt8JjLfsjr4+FeqdZnKZATAbPilUniHf
ar4teXlQzwvJ7fks7WzTtQ5WkfejKp0eLdO2IJgGdpOC08EbFsUJ3mx8T92155Bo
UENFz6IpeFbtvL91qwFX2nall68/LMy9hW8RArh/hBKYXXXUUufi2TLSEecdqDPp
Z/VpDcvU3GAxXkPkLghhEzGuGeI3zB6k1h0b0/dE1kaeAKZwsEr5o0GL/nQOOAyU
H0nskwc4dMryXbh6XmTr1UnyGRjg6tX2muCDvuE2A5SO8auHJjBA/c1n4O2oYhIM
4tyD23W60m/c+rJef8NtjfPJ6y/COMrS/boTjXM1NmyxxrxrlZ3iIcO5ZWroAYCe
9y5t5VvBx3t6PiYf/L9TWk39wXlh20O/WpWl/UZkNKMeRzAfCjUbTTksnHzpawZt
LmdnNwZ/Pvm72DPZJPgDvq7f4zxpdkdfxt3HadaPZALIddHEB6FnvZkqXTpObGQ1
FPFYe8nMHXgS9o4/V5pc2H8qT2CXBeVg4zEzlzSKQ1dIuZH8+DHGpXm9XRku2zDg
yUHUmiDIVgHGJLRxhCzpceY/yHWQfGwAnF7cmlhtdDj1yM/u21KCNeMlnnFT2UFo
tfuOXKfZha5j2UolpqX/3Ui8K0SYUkt0PJICGZdNpPZfq05EiOXZA44TlYjsWkKQ
cyGOWTSm4EgTbvhvpJ9wzG9mQ43H3WGBpYpOuppYR/i+2IxdI8y4xCuSAuTPjA8R
G/Xv6mNYpgZfAYH1ne9rok99d2VTJFATmJOhStf36I5pvwNlWmkEuUYBjfdaAtAq
HDumkiNpktGSjGD2YzOnyLDsP0hEVISgoEbLmCulV6pkNFDJZxYJ/bZiTS6T/3xK
S7lds9ODFQQTlLicmgn1n9REbhzS82XWMtoTUyxvXRoWSohqaxP4i/Z8AIihVW+1
XSj1R6S52vOdVfW+x7a3Pf6lNydgN75jmrLCh98QQDlj+zWxEKnTO1m4wI1n6eF/
31vWpergelZ/81BsZy3JwUK0GaatzSPNt1qG05JrXMbynIqC5wlAvmejKyNumZnL
XMgncNNSI3kFD5+1V/oqfOF0djmairnpsS6PndgB6fzstqNKk0YDgp4/00A8Zval
RFpsPazjMKqqN3e3O4YpoqVAyeQpwF8inoGd4AYNmYa0wEwa/lJalzP07gh1WXPK
uo6SpqxH7LhlYhTsbEFc75xV6AuGrDFG0q4014v2sGzD3JinxSDweROeqKwKwqCi
hIs7R98DoPoUzhhjNW8V0BKpvFuz8nOFz9boIMHNP5BYqFXPSsDeKBsXdcRmaGOV
Lil9tNyQ1JuU/oI2nLmv0KpPgzKaLo+Iwq3XBjqiK1rCFqShfRr3nYU0XjJcd1pF
cEGsUrcoy4fQONiApxR10BapoAs0CY+Avr60Zd8/zVgQULZSuERKB5uRY3zgMQLA
aXzbcu+R/Hww/EL7RzBXtlm38ynCoDdIKurWX5ViX3pdMLDQKpBJBIYJg8ZZVain
kvVjk6jzzya1HpP7epfegLk0FK6ZptvTLoIv+9xal4fnjhsR/dgoW9CGJTpSPQnU
f4rbNr1r40igrkxah++Nm/4ReVKXHEizj2sTa6h2LdtTfc8RjTqcZZscxd5T8Iqa
+bqL6srfoBh6G/zGKSV8qJ9gUPlmmDYKv6G6xIABR0ErCsNQSGI3x4tGveICBSOj
foIuUMiL8fup9E2fQp/7MOqVl5RQdRe5Gj7eM/i/TfjV//iAhZARxtFKtIeSS9Ff
SflEklzFD3eZPvoIsV7FA3jGnlI2W037uP3kc2ZV/VsOPbzO9gk7/PWHj+774psc
lJP1+fuLj+opPpXlG3VqSqbpcy6sfeF3Ad3abQruT6U7IlI0DPeSfRpIBp5x/xP4
W7g4BWsPQjGf8RRwwww6M3HRIm2ZNT6H3y16uf+4eIx+9LqpMcXGrlNU5clEc/sV
S+V5wKWOlenfie8MVW48hDq9+6B3Z5wtsWGkwDBkGHE4yF1cCQewG+3qWSCWryyb
dG3cgsdv+mVtGP9UzkJ0UIZSWe25C+QOo/ONqqFyLf6enQyTR9C3SHlYJj0vJL5v
hR08BqsW83zMYbfl1RbkFICrCS5DePIx/GBrYs2GjmWDA2o77hhBsYMTDcrReAKs
Nl0mpBbMm3fwoAobGaLIP3m4CtUZ1wuTb9xAasBXve1SteBSUbNdYkZM1ocIpcGb
b6zoa7SHKjXHDpY8Rt1zYFeHpxVgRfV5ruMagB5HsZ5fS74vpoxxn77TLUHA6lpo
b9TICvOsP9yPmQRzeEnz8f0A1SpC/jbqGD5hkr991S66U4nDsPLZrYI9cDdwo98p
gZBDgA7sTQBdfHSngqDm90GJcXYVkXXZKpnVZfWskkvpaMegHFZuH1uNYn/tYHKp
IULEoCCx3Q4inhfEjSC/p7XYlmje9mbr1PphJHiKBsNuyf30TXkaBQ7i77B9lzzV
//XHFfkV7qcroVP6XiPuOw57OIYV3MkY5IDqHyen667Y+bXjFFHY+2zzWlFfgfqD
yd4ld345/Bt7kxFwG7bMH3jj+27TAxG1JSy/U6W/fP+49hD+pvRLeq82+0shUzha
eDWLP0d3MDowvgMt2gma4XXL63TZ4xl2AheWQrKw/SruhZ5Q3MdVIbGLa5huRUEC
iJiii7X5UtodZTPv9pdxtOqteH34NYBhXTLNu3Vq30w411L1CpHRd34FbG4jmx40
8wQsceEuANTxUyQV056D7VPX6v9zJJk3Gu8oEzs3Jv5ZeTOwZQOJtsYzxKd7kLEs
kjM+MKp4qw/LG3ffXrX31LYTJKuyf4aJ0jiFH0ApDrl0DonN2MkhHjPLvGV0/3lC
FVtVGxmZdpvn969CDFfG39a5Ja1ToswK+0BM1yJKfvH+9LOStCAVgd4VqWgCHjqK
Yz52naeLdyf24UTTJX5e0oL9qCfLKa7f/+ldO99L+OnuRGA28NHM1mOvqFkDtnBL
MpWDLzJZ4HPQIySL8VAvNbWgoXwlC5RwpuKWYcnEg2cF0aloiowpJsCQYhv6zPME
ktoHDsK/inOOG0NFVe9+6lVTKabsCmk3W1G4Q308+rAaSyqo96OCQsmi4L8Lfrne
0sUNMfEB8C8lIKERYrr3oFmlb21kQv7BDa1uioVMlKw3ajO1dhKW4O0+TVRO0MSz
ktLb4evSyamQFqUVzFna9YYBDCGkSOzRNVhfJks2PDkMpN8kz0iZhIA1J1uVNuKS
sa2gRsjv26pX/FRC3o0nUtmfQ9AyRIq4AWX2FyIoi9AJ+oIV8IiNdbPSMnkhHfQS
TGFn5agqO58kZB8KR8Nlt7u6l+eyoRNDo+SIQ/PDZYQNjGChLU4xuWG22F5yVtpl
pr7kl/QcGhlX6Rhor3MC8m9L1fig+7tLPr8R9mB2IPSO+YUDDU+MeWrtp/g53pgz
zV+ID06UhdncPktyQNHUNQRjwGhbgQLxU/O/qh3ZqIZSwYMv3HdI1eG5TNP+6mc2
3Ix8eE3WAUupcpHb631JfSSjz5gokRnwp7i1alfqOeeegWHehpriVzoO3LZAkNWZ
BS+GRJg1E4ZKLr3fmOTX+qW80SvzhWXx8DhEFf9MF6LZDm3cuu5WCSisx592tFLJ
1FI29BqKR6ej/+T4TZYZByt5O8xM+1kmovEkQdQb1BW7mHmvnUDMSXLt4xk9MMlW
uv8QH4GPgqAZWs8kDugHu0yvnctM8F72RxNHA+10HFCcU/5wxRt1EuEyGbxR6JCb
kxbgqvVCjtb8cQ/1PJNrGn80PfDhw6qOcP/JHkt2U9ZOzzV0d6gj7vh2iaIZhTLU
iXkF1g1bLVHG7rwdraI/cs7VKjF21JrtpyQh2YV27RLixCXjDNx72XgM8jGmI0Mt
f6n7h2ufCvfaaEwlDMMja0RPDNFSM62XLFyTNyLjQNXs83IPJA9yZZbUs7jYckjD
dqb2e8UfWDsSW0qFTB3CSmolDLqEencD9234KI8wRd7mH6i3KpRuA00wEWStiNY8
r0YFro1JeqotTo2jDG8weRj92+03vfyF2Vca9z6sC12mVpATKBlGKg5tRg4ZooAB
W9oCmFPMLmFcvUQ99eI4LTbtmCauTI0XuDsvZO1iNgz/FFRH5VDfPdOKl1wn3qMN
AEU7v5zhTxLjrNze9xJMAULi3IV0qfaT1YxAQiUPMjIGe2t7aqB/UcOFmBA1ddOC
LI31IBiWxAhzaZoCkc/E6aoexYDF3P18vj0tSR9/9EntYY6yr05cbSAR3JluI5Q2
taexFMgTAaS/lCe5nHDgP+HFPA6hipY2r3vpexIosh7vFy4biKHBk4JcEEVzXoko
KqN4JZ1qx3zVQ88zrBUWzhNcyiW7BB7LgElseRNCSHphPTQ1VKOmEb9pG6nXAmFh
wz3uA96E8Rl1JNDszMi45UrWHgptE80cpYIj2Pl+3dniN8q4ipVdf1gN40mMJp9X
A08gPAU7cZSRwwcNJVgufta1Qd01bQoZzZlpXc+dFILRfy9SIVB2v2amNZVHCTy9
6GI9qjFl2ekbqE/J/uIQvXf24G9FR9U6f+fqCl0Lh1IlXn2eSlXyV9bGjCLdqmrF
sXnU46SpPmbl2gceOfkdg81gXUOIIyRiv4NDUzC3LET25KUiIUej5qawdb1Y7FFY
PqEJo6jxyJa/7XagOGQPs2f3TB1fp5SbJ2n6D+sSVQqPDnRtTOJ1Yn9fiA5Cmw12
3wtdxNbh6fwGRZ3AkJ7TDwrVFlSP4v/M1wHdXJifsgBZ6rlPeAERQ/Xd20+/hsI8
y3/po/AI8DXuR2UtIMk0y1P2YAqgbnPZKLKGb7S22w4WtY56e0qRT19W/Kt3uG79
LTQ2/ujIVgY7u7TUoGjaL+/O04fPCDfGKRPjtjlzTbiqris7XOd9Or3XoeKRnMO8
EnF2WF76aaLvg4md+OheqTf7kHBZcLc2yh/bkCjhWiVFVWRoAUHGWLM9pPsNVZlx
q5FmJKhb3rwdbHxiUO8hoU4jeklatqMnhE/sXEYobcFdXab4rrExFsGKx+Zi4Bzn
JDQpl4+xcP2havYbgQBmoZVgVGxsplAkP+Q31dfP7iKazpBGVCNyg2TCfKmqgrvz
iLmYNHmcPktRE0U9nk3Ac5HYSu4NzjAeaeLop3V77L6v1T8h4XX3DlJ6RQBTfVti
wO3fUVY0lqP5KSefaD0bT1K3OEGFhmmNSV4yymwtL2FdcSZow389164ro/nOzouD
8lcRlvcmIdoc7fI5v+W2eO8Npq6Nn8Fy6ncM345f9DXZ1t07E4bvkCd2UHiPGnou
sQTXOvbNxCI5whOBkolxIybv0TxAoiZNBZ/0LzMJJmWcp2JDZO0iJMFQsvfSslXj
x5Et/hgdKYsvwG7jl+wfeZ10MbWRA04bQ1t/1pIEqm72qvatUCc1bXh8myCevnSV
B/fhmuX7RzbhfvJECfZJTtwq63weOvIOIIwrOK7c7+XYchYbC7Ek3sQzfjBnPoY6
6qgwvaRfK7FS01E20DpuxJT3Wdk6Qpz+ov1wE9nw1Q199XHz3Z5K0hYbBbutmX7M
CYBLbO1gk8BM5zyDncrg3buX4U8lCiK8mwDODU9EmBMtFKqKOCprry/VYDq1bMJD
4Bcd0BTNAjwjgccKrqh4MVR4aEuk2E91lJJYrQrQMUbnZtzPtisbjfct9cZ0HUSK
jwcdrkoJ6qFwvF3SlxhJZT7FNhMku2B6mNq/G05Dzf5eePW4o5kQUT1dRvzXoB3Y
mo3ypmtjTaqVWeGd+nLfy0lVoCUHxWU5xfY5bfuw3/3+e5jrr8yACTGlWMnqzvtC
cRaZ/46oCVLOXiZZbIQOMKHX6R9yXn4x5+iMFU3Wd9brLEPrC/u+N0TWPrlrM1qC
Zuc06QUsY+Ueki2X/J95+Fr+yQNY7EZgN7cYirnh+dNv3EQtlQDUNVp2eGjh1qiI
xZ3DBF6n7r/TPcQSqmZr+/dRBpQ+nWhT8vfCQXH5JSU2d1IVR//xO30Bf4jN/Yev
NzcJmcG+xToGNpgUVCOExSQ4w9Kb4BhuxddkxVTRYuzN4RbGU777JmcUWVdD5LPc
MsoU3N6rumrxy1xiePpJi8NBl1OLYynKVHSSPt4RRcA2aXZzmmWpJsM+YnT3mA19
gjEFByYe047TxEWMEVoi1pVmq5KGnjuhkkvV0o6OGLOVWn3wDG+UZmCSe06ud24i
p7ssHCVL0SusRQFzQouRXhs0WBSk48taG9baTfCf3JDfIU69xmrjwyFtgztLCYXh
Ma5O69PRmsLWl6qIu8/+qkJ59+nsKhyLfyrZZW/DE2kDI0d3LntNCNGMZLqyuHfX
F5pis1JNpEMhX+IBm/Y7XsVf9vy82UpPfXB0KA4g5PDHyat+/+2pqbvwCvpLl/su
5SMtFYcze5Nr/IwblNgj5HGWaX8rdD5aQeN//Zr7sSMlP6TLxPlET+hrsqh9UkeT
iUz/PfHXgAWkmGfRNEG8fVAKcHP2/O31CsbxeAPCXUT6trBIF2+LorOxeKVzygwO
es/oEGw+wJG/AlD2xOHPKF4v6/SqrV17H6cIYAE0w9OtULFwhB+VwxSUc8jRGn7g
rt5Hwit2AFbr4kLs8+gH5a5ky1YK3N06+St0XW2KNilSJvw/WXAa6ZGik9+a8ca4
GoUqTz0Y0MFsXyxBol8YxI8nae+5Cjx/TYrLjTqweMC3etAyqII9tqkbyLgYysHk
LW352SV8mObs3i7wOfORiuR0ab6r+zibC6MNnPKx2qqAkL3dtQYpiv495XS0t7X8
X1vqIg+jXezq24P4/Dib6wYfG7wVPXlSM5cRrB6FD4ncis8pOHUfYY5YheyeyGi9
rV02eNlOXc0TDYHjvGbRPuLqN8h86OSl5gSlQTIgep+XKkwO0gOxAeMtPWN/UkaO
V/Bhfvjktg5QE+WP9KmqB2oEzT6TDhZ13yd0ygA6enxXuULJ0jGxzRrEj4RlRO4k
0hjjszazW6Joy3P3eyCKD7MExDY51VLByqLsPlfcMNG0xki+glIQcRJ3wfTg9O0n
sLUHBTBLAfM6K3oW5gl4aw9J90XOb4AFxqXi1yLF87gZp9pP1OcNlBgI/W9vDeE0
gZafHfWES3JgKDSXzzstat9QmZWe30RV0B2152DIVfnNh+2QXKiqPplqJ3PXedD0
YrNImsRYpYbPOOrOEaHBnDVQdyFVumnsn+9tE6mqLl2qpJPWSupqhRCKHgXohUS3
HJXKMVLudI4W3JHycdVVON1ZYJOZDmfW16NmDyM+sIlQKWsCfAv2qxNkI40vCoYu
enEw8wEhDIGjcQvBQqIJLRxWaGd7+p7MeMyMBgQZ/axWqHn8PXKolkGxF21Jc0VF
GE1Fte4pBSQ76QZXL7YMJ6aGrw6+kaUQkmXmkQO5JB8KfjCVemdbEaxOlqoEKpsf
Jm5rNNal0BK2Y7zHDhj9Nd7AVTJJtXfl+ecJxoBn0ytO3rM7dmqkCjSiFpBX9lRV
P6VLLkIQp7qH9qPaXx9xnHD/SWtZZVPcRvrPEdcT5Tu0HHifurXooOmlAvVpj4b6
v8qSWtrds3QV97jYAoXbzz4Fa0SNoyf4HB80KQXzVX28sNwPu37E0T1HynwvW1zm
KvKNdsM3tK+AVzL6A8ZJvg==
`pragma protect end_protected
