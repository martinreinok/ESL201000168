// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HYM55V(/OHFV?>)[6S\*X6<E(XH+^*OV"FD<=[F&5IKW(9+6]+IG8W   
H@"Z%R "ND,OR'FW<X3+)(W.]!"X'8$9=F@I]H5IFLF8P5U?4O[0I>   
H/_6.>4Z4DT'>=-))/*CEIS^QW94O>W)Z;#0I5R0*=G,^A<3<8[(:0@  
HN2>\]7*6-4V,S*P1] O+YHBY$25'IHY6>"+4TX?/]<-^<AUI-?PNK   
H $S3/3]MW<($H9R<SM[<YBO^$F8JCT \=>BOLE?N?3;1]@Y.%)SGE@  
`pragma protect encoding=(enctype="uuencode",bytes=24832       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@?9MU(/[W,>)U-5+4MY(O>=)$9[%K&FG?YL#@<!DC\14 
@9CNKJ1H!-H)4=Q_*\\P,6Q$7MV[(C3 --E$5RQ-$=@X 
@KEG*H,C!JS.HD](&RY>]0@G2P(]Z'"=Y*Z4:<Y%1JYT 
@K9^/5^N<YD_Z,K>:-=5$$?C5-U/\E1BM)=1LH<SFMZT 
@VCLP $5ECUO')Y8E4&1WYDXO VN^]IQD,K1E7(,A$'  
@:930BY"W7TQ>;R<*Q@VQR3@D96112LM?3<K('W7;[.T 
@ B#>C6U<>CX".,\F%X;J->2.]:5DV,?]OT8/$>;\2X  
@$V3-52=TT97$)C6V]$H1A3G._2P]5T?[MMEU-=&BTM4 
@,NHK<M@%HDFC($3FT-AOF7*US'5!V$AD;<'X%RF7_#8 
@/<F%=3CXYG84$NYOOS_2&!LSZGL%D$R*PD4?P=;KD84 
@=RIYU2+653HR. +S -^=+T9A6R[>XAET*'ZJP07ONLH 
@'=I>;%E)OM[8ND: R@@2]N9HA(H/Q3^!F^7R^/DT#F$ 
@F@2&7])JD) 7 _]#D'?*]8+>W_(4G@^##<N08J*$8#L 
@TBU. 3*T.3"T>:VEW#&S43;#Z9?PZJ#(._0\:VT%-D< 
@RM48+(*S-N1M80<+*:!IS5Y(S-O>_7ZV)G_'Z09]W&L 
@I>3'5_<&$EK7M28[:9@#+V01\0YJ@H_^YNI^'#( WM4 
@DK^'95&*DGRG6FE0A DOYY12KYSD+G/W0!?@:A]H=54 
@,N7AU,&V9$F8Q MAHG^  J+8*WR;S%Q*X+G.UPR=H1L 
@.3[]'L[#2_CC$?:8GF_S_N9\O"T&$+*QDD>I[6:JHOH 
@3$S"Y\GB.$006$C$ '25+:1]+A%&$)M:HX8QG'=\C1T 
@.[-O0&FYS4N1Y?P]%6XD/8W$C>H,\RDX3KL)G]3Y<Z< 
@[%F@X\,J0^QF<JIRV70/XUB!-'(7D?!6/Q52\;L\)$< 
@1<O/HPJWA/N!4F#TQ\,-O>T<*-H2+:SO/[1+"FT=]9P 
@)A3T4]X6!O7*P(P+<-K8S,9XL!:#J<> 8_K]ZO:TV_H 
@M*M ;NUA5G86@!8MO_C7&6$Y#N!:!8J/!N'%UL896_  
@^4 ,W2+AN4!P/S2;]4&?@DXZQXFCT#"9V>X#TA.T$ZL 
@^@[SOWEI/WA?#<Y4Y!EJV6C%A%W<RQO8?IL/H+#%HAL 
@(,E%BGW42I4_<4QA5B1ZGY7YYF3/UHF^^*0)?V:C@-\ 
@<#]%_BO"C!\O@RQ1F.E$M#/KX7 %HS1-;RC/8Z6\>[  
@L]"97Z!\5L%P,FSNZX<>\&KK[K1&OFEE;#6K"\2:B4\ 
@[A(PR LWH_4N'.B1FO9MB?=P*/5<?7@*,X6QM2[G ,( 
@(@KYH6H!81S/0#=+J33?SGI9%Q=F">:HV4P%PW]CT_H 
@4G2JZ0%TW%IVO4?2\81< I<GJ*#P"72:3*\<YF0BVPT 
@>AA\7W[K#(78@6_C/!U[)ZYV!=?Y T$H%H&I![<WB-0 
@B4GN;RC$7F31P8C6K^6"4IB@8TU+CX-'JO]@9+8JGN, 
@W?8Q^L1O=QP%=6F#O[--^'];-JDL["];"[/9CXL^<6T 
@CGV5TM_SV5L<?)!.NTGDOX(3M5\QR<K.J$9#[D&F@^X 
@4K<B6?D$FH$EE!XA@*C<CT7/5I_@Z=X1JXD]9U&"V%T 
@6"@W>*J;&5!>U=X>@EAA7!"B;7+8[#@:B(MIKN;I\@, 
@L7QFY(M@EIU8H\QY*0*KA*>"2W#A'E<#9A=TN BZ6WT 
@4QQC*19#8+R_T'*^,;1_8E2_]9=2Q$6\(N2-E#2L,\( 
@4\FI]C+NE"5G67_@H5EK[)BV(_60^8V/7L#F6RX-J60 
@#],:8>:S0C603]:.V?,&((\^X[@P5K;V([/5I)>\$#4 
@OC! P"HNJU0RQ'3] >#Y6_7<W?XX4&>9$E.36!RO\&0 
@!N(A/AJ-@'V!$,K)&O_*L[<5K^[+ @';.5_=6#=&F0X 
@'5?WT%$=P%'OD1?UJ;?I+W1O_Q"\SW >U($!TF?FIZL 
@L_7_&%UY[@777T'0^T$495[>&+W SX.=4(F@YM_-07T 
@=;?&$$Z77\_PI.]T</3YJP<7L[M#P HE>W3E"/K,>-, 
@=@*!9@CJ2UCN/6^U8M0RX]D$%!2B5S2"BLAV1UT&(:0 
@5L04WC!IJ)!^M\" ]H3$'#@1$EYH^"2EJ"%N<=AI^U\ 
@N0VKF@EDWO<7% -R!1- /KKO<2 #PB],(AO=7+Q1)C0 
@-@06F!RXH; F>8[!_8B2G4YNJ94C/ &Z[,YOYAY5O:4 
@&:E>OE GO423;[E*!3/O'"!H#QG@L><OZ5"R10LS#ET 
@7#B](S[MOVP3OJCC__"S0UR0=%3:R0^--4G-0NYS7$P 
@S:?X!"BM!Y4=TAN7J%-5Z\^"7H._7F*X=HF% \4@6LD 
@@%)&)2 .7HKJZRM"5C^)G,,1E^9AOL_"[E^UGR-+$*@ 
@[K&^GE]X'#-1_=KBO.H=G]^B3XBK/&+NY55FI$, SI, 
@*$Z&][5HU7YFP-(OS!]E#(+F6:5P! ,/?U&M?FPE6+0 
@[V]_:M+0L7ND]]!SK($E)G3F-M#7-2))4K5/'_UM>U0 
@RNDKX6FQ.54PP59T%'F;W2)$HP^DV90I*>_(UB_ !-\ 
@._>7J2V&%OPV@(,3>X0D_LFWJ"#<HJ@BCDA:CP[C2JH 
@ISED7*!?4HLCXHK%64\:>RRQ?S+Q_"R9_H:>JYKPGWP 
@X;]WIBNEQ-18*88JAMHY*Q/4CD=J-1H]6-P^!V+/D_L 
@P9D),R-DN0 2YS?V7"]!T0Z<Y_M*OE$6(-6]VQ-2ZDL 
@";Z0L0W$(,W),=!24?S/YEY%A:]%$JYZ^M$HXJA;W6T 
@AHW@@07#]4T^P&TQPNG $4%0E% CH",=ZVJ_71H6H54 
@7,-J@EVO%N\&Z/7JTS[>G)[H!'10**;KBT_'>@S+&N@ 
@=>!1MX@*NN[)'^*+@W1>1W W+].'XP8^%!L>.=9*%#X 
@CW:L"Z.6<H9K39U29<9"223(4MSC'D(F.)AT%!+3*]H 
@@KEM%13P ZA: "MR6R(BX^^_ AD4 6+!>N>,AVS-I>X 
@93!'>D:9O$N:"!?6>"!PAJARI!M<BS%)\E.AJMMPQ^, 
@Z>C<.UEG== =HT#EHUVJ7A*D[,@HS1!LFL((A @Y FX 
@R]F-48]XUNZ4\'A1/2=-9Q_A1%ECY%C<C;EGJV,$ZBL 
@@T3R5P3F[=D?-V\'_8].(8"^#[)E2$MQQ(<!FLHXE*T 
@Q@D#,7<@1J2+O+FA850_:>V)26M5&W6<+ ^#WMY&R0$ 
@\.AET2J?[*[)X6YJ-Y^]KNDGLV#[#4-$ SK$PJH 5CP 
@J>S=?IA_]MIZ$,SV8[[ %=):X6-EH!:L<>V*$K -4H8 
@Q0MP<< 9)'XV#B1TMX)%M] W<I@SW9MK]#NE:(90LH< 
@7X'E4'#7O[,#KL)QTA!WW\>TS<,_;?.R6;_UQ<1G$1\ 
@S.S_*CE9W4U5UE$W"<@^,:*X11U&!17-12%L_3<XYGX 
@M;JHD]3SL)K 31VVP.JE>Y[91&#V?6L*18A'L&^\/WP 
@>#+7.L )9HKB3G"S/%T4X4?7_F$^J8<9[+_2HEZMQL\ 
@FX2\E<\Z".?]Z#)1M!&;J0$)U5& >ZW#)=Z)Q\'5S!L 
@GS6M:%U;%,F-.LX_4\2^1&9Y/#,6=Y''%/&X(4"MCH0 
@],<;TJ;$]-L>:(5.JV+ADXTI X+LSB5$R;SZ12]I#1D 
@4B+WW:,,*'9VO8'X D<-6+BL!S2Z^629'(00R@AMCJH 
@65Y<&<@-:.'1T*OD[:E7#3>0Y_'@HTNODJ-+7-7OJ=8 
@T N?Z\+:SW>*!'2\:":73:AVBS=0(7XU$%Q3HDXU#:X 
@3IEXLE"#9THT;HN[,LJLM[DFFI@RX\(!4F26F:1;6"H 
@60*Q9FI@@L?3'['M7 %OH&W+1?HF]2JI<G!7:6/<36\ 
@!B:W8&H46/PR2-L\ZXU-AO'#T!11;?.>^_?-@7ZE=O( 
@*F]"CGD;$".'^#UNBOR#"B]'\%&A68P3 0/A-C8KJ#$ 
@X1#4T&XR1>C^8$QMN&N4-5"&>UPRSP)+SO+W;XCI.%D 
@:#A^'(1/=HGP*2F-1/H9 E(P%;J)H"!4C<.OZ.0MJK4 
@RL@5WNVEQ/*85T!&M%;-::S1"22^])H\(75>O=*G3(H 
@O%\M[S-F/?9&.O6MOK_M0(?,N862%9HA_++>QD!F*2$ 
@BG:AQPG;L[C.9N-XU/K9KVSK-[H:E8L#MX!UI1<10B4 
@4L<NS)C+%;4Z0++16VO62UU$UB8<=8(:^%;EH!%T$XL 
@8J95GCDQ+->W.E\KPY'P=5DP0F@JMRNF//MM3:57D#\ 
@\S;7U++Q=+VB8"TA]Z\2^$S/GOK89]>:W':?9 E) K8 
@R#ES\N@?^)N@<HROW^IE57:I)%^#Y@_TXW#2.&@Z:MH 
@%&2%/JHL1$(\T+P:)+:BH&F4HJZQ2:",/EG0''/])8@ 
@]#39!S:7&VV NZ3/_D&-!HBA2K0]D4031+^ZO-)+'OH 
@IT$5^R"6B*0S=@_(84HE0M64?['H5!I*=.SE,PEJ MT 
@S#\C31T!A*0K?28I;.RWX;;ZN(O3^HZGX6&Q6I7#^IL 
@3/WE\K$W&4-Y0_Y12E',?1$Z03#=/@J2@=I]5D\6(Q\ 
@2'<=-/BA6>W"@6,#&,"*B@ ]LPY[ZID2#X)S3,N.@>< 
@JU^/*F?43,I>^>&>3C,J#5Z8@A(1/BUS93)U8WY$I]$ 
@.V*TGK?F)^FQ:YKT,VXYE=?)!8\MFA/;;,MKQTX\,AT 
@DY7U=\"3?=T@'&E ,13/=(R<P\PU5K&S:N)ZV6P!N)@ 
@0"N=Q2 ?Z]!MP2#I=/79TX$@@TBI7_;!A3+TZ=[C.Y0 
@@(2V48R3/0-:4#B-;?W=L+C"<RW^&I8EB9MS;[9E7^0 
@<$Y1\IP ':SSJ?;DX7!&"HP=E+\%_01TH2*5C%>&'?, 
@PWG(T584F'NB8<EF4*U&W3RN^01L<X]GGU/L"76A;*< 
@>0I^3NZ!=NON906HKJAFLC2H2%6F[)3#X"L"9?I$8*4 
@F>B]Q8WQ.OYAQLGF7]"3DI*W1FCV\C?'+?X<I._7_OX 
@T)7,"V#U0<W92 *(.Y]['@AX#@1?2U@AQ@<0M9M%R4X 
@-HA*LQPX<E\)C#*;@LTZN.QKI(,-4]E4K%N+M3N8\,\ 
@5HE)SX*E_?]_BMW8YF4 VBIF%1OP$MI<HFY1.* Z>OH 
@TF"E8*QE9RRWP-/.GF3@.J9Y+A"FJ5I7WR%Y[GDDJSX 
@8IS\C*S39_<J_U$,-> U"B,72IG%N[-W9WJNLQT'W+@ 
@?A0,FA5B\_$.Y^S4/'-1 KZ'X5(#[L_R?80HJV<50(  
@SVB4GH[X-H:3.B6CBTAL7D<9.K>>$AX26P0*+KW6B]  
@Z3)1VFO+9#E7" F\&*:NK0@G8P)&W.7X?:RZ+<MU-DD 
@UA7KY.]ED)+R(%:=H05PO9J\!7=!+5Y0U6T(&4<D?%@ 
@5[EEHD%-<VQ,GDQ! SF\09^;D)"M1?+<M\Q.!L CD4  
@.$R!4C"'ZN9R(4'?H0#ZYD]8PV $GQ8665# KQ4(&64 
@,X4O"=75B@,XOD7?>XP!KG5^IV15[SOGYC-BQ5]G<6  
@'SQ8T'A^?#X\6J7C1V=6](F8D@VUQ2R1.29$?+/S;;$ 
@25[_J^73]TL5PO[$QTA?'<;*CE)%3*L7&=F67.*&V^X 
@/AC798*:J5J2]I7B6Y'.D\P6'"4R*/;DK ;>%"@2W:0 
@'[17Q_V[3S4"AC+B\I8*[_V!3&5DP\@D) "!!;I -T8 
@)=13=F+3V[N*=_YU:O.>82ID8RX;)8LP<DYM;1WRR:X 
@7>A%M<77N5,_*\4@'EGR[&MSFR8AHLM*17TPQ6*^LC  
@AV0*3PQ_]&;^2YD_Q>?@G<5<R*F5-R*,@Q$);)4S/M, 
@.F$I3THA9TVF@&2M?U]1C;_PPS(. >@!PU"(>V^U=-X 
@SX9H6::IQ"9+[O<M 41;@/F!(N9FQ6BX>(IY8V[M"]D 
@^*W.N'W!S<"D=)V=HE:,$JK.7FG/96 $OS[=C[%A#JX 
@YA"SY%/Q(IE^!RXCFK;(0:H+57W[P3T[;^,;^0R#[%\ 
@/I5.-:"T6<]<0#$;J($#!CY?OH*L@% 6\+_ [@4.#H8 
@MURL!" ,M!DDP231GQ%9(M4J:\\BOFQVF#Y)52-GUAP 
@_H^.;2QYH*;P:W"]RC6ILM>GQ34CI^>X$O_A#_K4_%8 
@8:Q5H23"4$X/MGVQ5S%?WCJ#\G*/._6,81MO-[/@&4L 
@)TFF 1?N08+O8<JBH(\(?]E1:Y!^_Y#5K6JBB  L&Y\ 
@E/!6<N='<W(7ISJFQ>QHEH!S9G]]HR'A<_3#X@3M"4T 
@_F*%9^Y9:4AAHA"/>Q<1E9[G!X@.9:UD.$77#7<%TFL 
@_8\FW%>&!:==:3<]NT6+S#A,#DAK5=\LT]L%H-<'SBT 
@3-E(?T)H7?MS.J$!W0UT1NO7!K@)1$8=(7ALWMNIMC( 
@8EO?1W+#U/,J"3/Y2/+U\DA0KBD TG:V6,6KEC_@A^< 
@,\VAX1Y\+8TRE)C$@]N+G;:<>RXBQ_)HV4S!KI596 $ 
@CL<-IU\&1X4)\32P$=_I.;^B09EY*;A9%9K]T2O3*#< 
@XUL%! 6?>_$$?PT//'&*1' ,SJ@0DQ\WTJ;1DV68S=P 
@43\)$8&2-CJ9H*5;7Y,Y@U6FLR(4S 2I)AI\130TNNP 
@J)^@S*!XY'>]+O(05OTT#5I#J@CF71TDV?#0J0%,-P, 
@@O#3O[<+%A5;\]P1[B6N+0T0=)0E7,#F/+94M_CXI^D 
@;T9;O;L!K(LIDK2J_X"B\H?.E!M$!M!72?X3=EV#=&P 
@!J#>=+$X[M:\CWP_='"MG_KHU64Q5X:^>\;8.1B,X_T 
@:4<VLM++#K,X1T:'B;>ZD@KVT,JC?3XB<S[[EOX &64 
@*['_=M$7&P@N^4V=4PZ:D$W4YOC*3T5A:%U+C\@4Y60 
@59B7,'9;-@(AJ"1XO], K']*^Z+0'''$V M?S^;F9RX 
@#&".EGV+BU4TI0NNSZB<YB2ZUM</NU9WD'"Q3=-0'3X 
@S[ZE@U15"U2'!&SR8+/W.1T+<H;.?89Y9]-&DW:,N3@ 
@6LQC@0MI)+VYSB1]ZD7DMYT!+\%B'8C7F7Q.,E)ON60 
@^OBF7JV2BQMAA_]Z7)@?X/*N]2\.M,4,%K+:B2%Q":0 
@$8HRH1&)QUW;'U$4'$4>)2# *R*%9(271]?!-;P8Y>H 
@ #(]./3\8)FK^\^WR*),AYM@?=DI!W='[I0#E^DR)1@ 
@'*'7J,BGD/JC-+Z8*T/U'HB7'>J?/-*LWV)\GM44"Y( 
@C2AP]B7I\O5[\BM#!4^:Q=P]588N!XP;ER.B Y/92]D 
@[M;K$=,K2^-2\N$=34Z"P;3\W'2,X>!*UN;F&$6?GR\ 
@+G&3.)41K=K^ 2-^,[]@D:\;5-P#AEJ<SR;E\Q83K'0 
@P25H3_\F-CO/@SD;7*/5.V&#9(;.:M^ZAR+HL>_6%V0 
@HN^L]Q)E139&"#RP'9!0:S6% 93+0K@VIB_1437D;)@ 
@QJ"W\C&.J+6,@)F/S);8T3#VGI9('C@G6$''H(-<)1, 
@8+,B(O.Q%Q0=#3]^M4=,)'[&J>PK1R?7FYF\S$Y*!^( 
@B"=<]NE)/"O7.F9RT>U4! -0#DQ]#'1JG1S '(?#HT< 
@YM0 */Z*T!%C/F.*E;5J#S*C.BNGY*TB_M>%>I3N%CL 
@J$XO#2^ #RH()(!F_\^Q/[=RVSJ5I*VS]L U[@6'-U@ 
@O^#O>CQM_P17R]4Y)B4 ,$2*>J$&O@GD%!*/^@E8&9T 
@Z*+W_LW"*T+^38IO8BV9/*FZPCE8;.KH,!8/W3E9\%, 
@T,0$B ;BAIM^F.=\'%Z)BU'BKT[T<3NV<1A2Y.9H75P 
@C?P)+,#$5*'0-%U$H2'%\63]Y5QG9OXGVA%<]WR/<)T 
@>K2]8IWJP+ #KX&+MOV6E*:V7.#,P:^%NX[-LQ5A+$@ 
@JU?JE\3_NY<1N:WI),'3*=8LBF1EEP$:/:;UKB$7GAP 
@:[^?,UFC@I85*6D'"5TS:M/&HG]V(D!KMSC.@8^5U&  
@>9O0N5KD3HB1PU7@'KKS[4=3CYK"ZCFIY-#;_:#:GND 
@J)MF>Z"FS,UQ5?T >1A0<;]9-G$9IAJT;>LI%B;3=(H 
@1T+D-50Z)8O7WRH=J:?ZNJWNB7]PG*_)D5O >?Y$N3, 
@\8@A3UI()B00U=L",.$9!C&^@B4=F+6J8D)LNJS^]9( 
@_O'8?DT&OLYR\:K/(O$P7AB9[@#"VR'EO4T_]/-^.H@ 
@;+<<Q8%O5:/"\#4S%X.LYKY@CSE(#6B7&)EIU[]+BJ< 
@;E@E$=:_)OFCU=^$I=F8XEDO5!4GDD'XBSQMM9^#QD( 
@R.U)TZ<+QK>&T((.R!0N&B@[V8(LW!MBDRPJ>24O67@ 
@U&-*'>R_G!ZT6#8280,M$IR<,WP<:+!0/S+L%61_EE( 
@K:+,++YAX%X6>^%_FC< M?BSGNMII7Q]D G[R_M)XE  
@5B[N^T(4(Z0Q49\RI; $ K9CL$;WMYH-$&J;RK7%#K< 
@5%N+(-%"@4(,CXTHXTA+$A!L0SB&A%,P"SN'^HU?9(P 
@^*F%7HNNIK^BR]>#)^[U>P-MWG2_V[T3660 *N?0_5@ 
@>#!BC,MLW![LL A.9M5N"V>40Q:N2:.W6\/XQJ*+)#H 
@>); 3U[2"4QFC.%0>D+P:-D6(9<JU7EUAK3VY >!6<X 
@EG\YZ=?QU/,&7VR$:.:$4:*"H0URM5(,1C(=U^6(*Q@ 
@**3T9JM8%X[5"6JE<IO(MUZC/.< @^4!>$93!<C%LRX 
@3904%+$Y_%W,4AQWU7LI*WY(HQI9<:"R@9M;!%$O/\$ 
@:+(;SZU&,<7,;S8'*TDP&ZBPAG;@$1Y<@=AXHE6X;>D 
@1[\&Y$0S@91E)L6H5 F@9_0[LECL*.2MXX"2E/SYLHL 
@=2'I<ZYQ:.?HT0D9=8*:6!>S7S_&C.R#DWR3+-*2CU\ 
@.5YV0_@?=M)\)K9LU*)J M:+6X],*<'",%%U(X1TI@H 
@LG@F2PXLW]%Q7?\B [VB1PCA,"?<"H<7<#7HH!CN:=L 
@K8ACH&5BP0[J4(N8-E/>/L]J:C<>%R;2Y+QZ>V>DACL 
@5 NPW2S@/]K Q!NL>[J!^ZW5)1MH8T'GJX["Q>%.\Z< 
@EQUW";>JV\W"<VF+?T2E+*91<T1N007E2TB&Z!SL0U8 
@COF3J>4XX;II+I?U$1H>XE4"[;N%LFA',];F-M$_A.\ 
@2: /$1?K;R'F0@.VUBH-E>R:W]RKPYC[&L%X[(7>1"T 
@!P)1/=A]C3]C'VA;9CH3,L20A29H:'DKUA,RTT(R_!D 
@&=@/&Z R;L0M8Y"=G\;2=C=WA==P^_ <YIP@ VRD<M8 
@;)RZ'E+9@5)>,O M-06HB#I42.9Q0,%!ONO[P2)>WQL 
@BV>ETUX:>0B/34P:0-P9JI(9B\^CL1",ZAET).8=A7P 
@2N6<8"*="%\O15D[0+X\.-$J"205O,ZPGU S#*!X0 X 
@*EITL<Z3WK"9\,,Q92V?Q_JF/0G"D.SC&_C&LDG@4L0 
@02.J=>V1Y8;>!('(H>S ^ *3O2:0$KU(/S^B!MMGT+@ 
@U8:A=EK%@C.K12'U>V"0.:PX\4D ^QJH.DXZD!LNWO4 
@+BW8P'DY)!4I5ILS5C$Q5)!Q"J]R CSA%D,_$IMRFM, 
@]&H!/[+U J-H,PJU] $6<)C-9PD ,B#7<D[-8V31!;@ 
@$]N?[NXD-5-[OT$L.NIN^E1WK#WZ-DF 48E?PFJ\[JH 
@(L,A$3^Z/%S-8!@<P\OT?TC)RMVBHE^50O,-3*;M7U$ 
@1U2&:JAE])!!,^9*[O<4 LM\?>SL0L8M,U6Y@8N7Q-< 
@A@3H1,G!T(IH ,*_ELL&CB0Y28?*/\H]&#0+A)$K\/@ 
@^OG[3_RLV!Y]3G+CTTUB1(R@6"-7TX>A@V)/G/K_K1  
@GCQ_#"ACARBM=03"K"N(6GA_=31<+:A>\FCJB,90H=@ 
@&=?A=ND7;6F1#6:%&G);M>&]0AHUAIN_*!!% =5J?D0 
@6G'L^7*[F'A<N<HRZWYA)=N[4C5<0G620B;]T^)G=GH 
@,NIJL5VCIID*)KXFA*XRSA49<9"K^?TDL!&>U,I].@  
@'Q_A>?\JGJZ@ML*+FEQ5"^$4CP$IJ8[?;/DJN&A#PND 
@I52C+^?VIVH0F&E+Z/1;E$;CPY5MNA%DD%(M3^B3,%0 
@B06332CB9<'5"Z7:MVM^Z.<NV;7GZ0\8(:E".O ;4'P 
@=C'N6S=BCON:!D-I[K3LAH-(AF21I5VF&0+"OB/7[)T 
@NXXGW'>TRC@_L"; PY-UHW[=.?1AB#=&@!=<8\?Y'XP 
@)>2&(X9<+F6/@&^R\<I3RF7'Z+W;#OD,]]WDA?C- >X 
@8^OF)2Z='PR\<L0);7729"8_(/BY&SN[0"@OW]<4#;( 
@OC>VQIY]F(,-Y_H0,.V&K>9AV0HC].UHRF^B@Y,PDWH 
@2HJ*5U\ !0TY)E#? [,?"'^RPBE)1S7*X):E<&#,F[< 
@>FF.]_K"N%VFSA$+PJ=!NRO=0C?^2W. _R=-L!/=R*8 
@C,C=8;<[UT1!.OJ^C!A%D!/%A=AN_Q2] +^YHD0$SXL 
@,2.*RC/PFYIL7SQ.N8$D#AWE+]RO?:LM/=T,U31E_0H 
@%DW""'LS\TRD#H5&R\I>,+$=ZTSXK&YICVY\>N>T@(X 
@"-%K9<)T,<E%)WH;EPQQ3GF#(J.D1V8L=@#&>#.!IS\ 
@"F+0='<=1 ^J\!"!,( -T;&U7-G;$3RWB3-7C\[0;[0 
@XA1NK8IL%#)I*M+9G^X,5Z09IG2 SYZH9&<4"=MZ"Z4 
@=[4R\K7^/DIK^4%=>>2<M1?1-R3FD->\.&F8*L5&7Y4 
@W;>DR3@TQU@T26+'Q_*;Z;]6=W-A/Z3.F:H4TD^ -R8 
@B+(QE)$JI+'9'LQ94*L^4WL]',*8CS/(*LYO1%[>EYL 
@FU]48-@[O!?/<ZV)O[$BF>2W(ZZ#$O0@J!R3-Q%#^N0 
@F:!,;:IKFZDB+4I98^'-"7FG[RJB&I-X8\SV#%\*L>8 
@O"(ES1$VB!\&\$6AUF87.VS=3R'LD U^"<' ;F#"X3P 
@4<WY/*/E7QXX&%+#HGSD<P"!]5U^ ZP%"92:#,PL6=( 
@54G)/S.?CD;Y=:I7IXZU\7<@.@I@;7_UU\^'3P+YI=< 
@^*\(OZ;+TAS]FBYX%7X)-I?1X'.D7$%/\JF]HX*2?X, 
@>M+S,8-;G8( L]*$FB5G!H*F$F @NS6ELC:)C2O/%E8 
@^'!G>HPJ3Z1R;:"JL=/4,%IVQ2"XEZPAP&#\D@35SQ0 
@W,JYP+3#7$X\)WTFSAC[J!.KRI+?  O<3<"A"C5?S]@ 
@",=EL0!: /XS=.,-AM$6+XG>4-7QZ3K.VS^9Q*RJ(8T 
@[H*'?EYE.6O+?%#JSS$2J$O3!US*@'2>B-C2ALQ>H!T 
@79GK=>&\AYT1W!H$OR0^]JN'EZ0&Z<Y_C_?5$1]WC_\ 
@C(> D.AD%?IMS=#.H2=^B@ZCB])BBH*82OLBOXGN^[$ 
@"^JW^@(T?+6JV3(."%P55<U&%J_LA6'H[U3/55JO5H\ 
@ODGF)HP@W1446S7-1..E8XPDUGVB$C.9%J,,6WZ8K2< 
@E/TTAF384S-87=7/R_**)8J(:07O@OG)3H16G9YG,U8 
@]4Z L6=)P?D)SV'I>J&@E PJSU9C)QRU%H6G,2 B]:, 
@C,AL#+HMXR:<F<J*]9E%7@IN6G:FP'N!BUPI/F;#'6, 
@\AI@\$#!@MU)9)4M*"1-GR6-)E]\P48 *A%+AI3Z<#0 
@1"R5"KYCR'",W-#W3.M6@@MB"T)EJ29A1)V;+"(#ZMH 
@D]UAKN38D+J'\V>2Y]0Q_Y\6[2+PKCV2E@\VBT4F?!H 
@!*=2*%)C>QZ_SF M ;U1KM,)^S/1)CWX(!<W]V(D S8 
@JKE*L/> 5=C*N.P-R+B%!5;7^J<]Y9=263J@8=J76MD 
@!-#0&6B\R?U!N3FA'\71A#91>QW>--@=I<502&!&CV  
@'1M4JAH:&CE:%".NUE%:4L>J?"3G"80<Z)[R!O[AW%$ 
@DM];*"Q]1\"NKY7;-C7S0G*S*4V!LQGR4_1OUVQO'7@ 
@<!1IL-=4>"1QO<(8)]N!;8ED<$/U?U&$84+:-VMF,Q\ 
@^AQHCO(H-<#+CC7G 7 8R%_OYK94)XJ#F9TFR#:HM'X 
@+^S8*SI-VWSO;0^Z#+M<$^JT;V_Z&RT)&S/ZC-Q\GS\ 
@@%F,P=P;9IUMQV28$,#!(6P]>;'A2VEY7.MJHHJP,90 
@-KX28Z%RD/#P#W#I2N$(*5-1ZU+ZS/12U)\3L:KZ/0T 
@/J]8AKZ#0D,:BUX\,0LC0TS=5I:S@7U.KD7GN]ON'%H 
@GMOWTH)!U\FF)H69&[BTMVX<B2]^M%7/6=[1XY -OFL 
@J6]*#8^I?&:V837&PMS?_/C=BL,\]4@"E<.@1[%'<", 
@JHU*@Z!^0[*H D^A6PVI@B;%CB5GICI(%O,W]S:%<0  
@D3SKJ)3A.?S>%E&A\@20]I"'3-@@.7)6UF)?_SI'2]  
@.Q8##*:!SBXLAI!KUQ3P.GPKNC?5%$@E@"X1I)OM>BL 
@N&$2DW().Y%HYDFRT;0?WS3 U5CD,3:4S-QFX+'MQ[T 
@/H9\[>14OMYAK,.^L&?#!T$=X))1>+2&QV"Y.G-("5P 
@NXLGPMIB87W[ZF'$@P"IE%R1,L(U201FW:N3418$,.\ 
@\]T]J/$/^\C#(?A],P\;_$L&M(]P2K&H>.Q[6'/K*>X 
@MR?##D=V_#8<1'."NM^H''+<DD&5L2.QBY<C^GPEE,0 
@(9 #X",L"V]W@!Y !\=K"=@/^2WEXC3CQ J\%*N5CXD 
@.^TWY^^^IU0Q=Y88,MFLVVH]@N!BD2CY3="@6*Z:"!H 
@$4H[U;@&(%$'&IYA@&B?L#-S=0]2K;W8]9K<3M3KYX< 
@TW[8"!;D N185GN(*$4KP)V&H'6;^0VTN:%Z,DMZ/ 0 
@P\^M=YG=Z2?V393C(T0&AV0 7JS."Q]]FE)+*]CJ_&( 
@UQ_T)AP%H9H3L-=KIKAL#G*'F5*16:5P')2ZY[#6X=H 
@2?+5!VGRZG>5X8DB^!Z%#N_[.\&%NOAN,-68&[X3>N4 
@IQT8H-65,\_>&>BIU3@/O^*\1Y#=I"\[ 9-RN1%[0QH 
@V@/MGCSF 7Q1!4S+DI[T^"";H>=4)W=FF"(W#5NC4_  
@'!.I>$D0.',3J#2@;Z+8Z$W.BS]:JENO7H7U]!N2BA@ 
@AW?:4*^)YTO8STES*S#M1GTA>;H.!1"RM&4H,;[!.], 
@5&HY5!I;X2K96\F+ ^9/V>&]X:"-3/L-G "C<E+)G-P 
@E"V[X] X9'$:4'9W5O/+QKJ^P@V[_<5FBWBS(UUWP<  
@&T+<KFZFQ):.XN%FZA W#J$&4TNP[?)JB=HF@E8^6[P 
@V34\PNJ.R1I2*4@JF("^3X.KKI1#+WDY\WFP:II*;$\ 
@5=>_'K:_AW=5XV-%GDY.490'^-:;$J[KQ==W8AMQK0H 
@CBD@5K?')^]YG*PF0WX$G#*#Z7JD[(&M1:(RI].K)M0 
@9;9!0?$D7(?2E:=_62FF$8;MIWP>:QIT9]$"7[59EHL 
@?GZK\&DS3? 37@2UB5GF&;TNM#8&-2+,B'V;W=+JQW, 
@YPT-/>%KRFI_DQO4+G(2J3((.2^J1,PIY4"F])7E8^L 
@D9XAQ]5P/?2<_8Y%68$( ;]N(0R]C[F@ZN=W;%X:T<< 
@3QZ20AJ$AS*MU@35NJ<WILW,F7,M]M")V3@-N;PKP34 
@^_["<00^T@RY-1#OP3W;GE,YN/MBL(S<' :J&L7N2GP 
@(^D(P_5"@41]=:ZH3O9Z8/#Y'>A Y**)]2I!-[:'U;@ 
@%)1@I/".M2019D R^7$YPEH0A5AR]YJ#W:!F)>P36[\ 
@.N#>COSX[<06I##Q[MNP5*H[?7S1.;CD:,S3]L#)J<< 
@L6>)7G&8 GM2%\0X\.:0PNKBJ6!"GY"7!EGWJ>A81[T 
@S6?Y?A$]*[L[$+(_NU0J'Y8$03:97-1!*UNG[51763( 
@1^!.ZZ?>5!)K'UWQL]2Y5!7,=-J< [EH]NIT7<2&^-D 
@3G9!DV*RC>[C+(-PBC>4']=0(,G[G!C-'SSVI[12]G@ 
@3\; #L[_*/*UI;=^62PH1U!=@[.U$8WN^DH2-H 5-+0 
@5^'$*W3$"LVWRUSKMRM5OT-.",^9?S[@L.O:L<U 7[4 
@,($VO=.LSDMB#;NSC(<2L"I1R17B!986%'AD?][L)/P 
@64&W=N2S[7[2RZ$DQ#:NAN++%A*04K<(XTF[BI:I)OD 
@OS%0(]EHQ1AR=Q6\ B:>@/Y4&.J27MX"&ZQ5'ZVPE\< 
@XA\]A(Q2[D& W,XH?AG3NK?[B'4"Y272*<NN?U?.5+L 
@;>3OTQIX48 SF'FK*"*6[[D")H/V)@?*T^3X I?G5'X 
@'H G<1H,I^Y*JUO0]I''?V_^@13/#3[IS(!(O]0=Z!$ 
@#0+5HXL/7JD&/: \SNG$B&-*S,JD!G: JOZS@A5-=U< 
@F5OT3RJ#ZY\=NOF5NGVXY<Z,ME;3AN,4<9'AD:);R24 
@YV)'N$VX<"Q8#+5I_7OD#]>L@?S1L#)"I7NM#=),7)P 
@M7G9.EZ/J(;T0P</IP<W\<Q)O@%RX@)$AII11G34QL@ 
@3'"VC&5?RS5LZ7[:5:^8\E[<]ITAP*[]NQ:XTKP3.5D 
@6KB* OZ3=R):G;D8 ?]"_=OUBP=(1Q,^TQYN;DL$UZ< 
@X\W:WC1M/]:*]9GFV$, "?CB*'=K=9*?8$RG/4VU3(L 
@LCJ";H=3JQ7KJX)*FFW2X@)<ZS/>%FS>'';$3!;*TR4 
@+>^CV%<>5J/2TBHCD!J%%ACSTBPH?&I?PE(8LW#V,'D 
@?NKDWI@]T.\H"K2?6_"Z+J7GL=#& VH_^R:ZVX[_VT$ 
@M[2!1B]W7'0A@Q%^W]C'GN.V,ND$DID;>AU>$G'^<KT 
@YQIB3$4XE;+43"-;<<5)VPOMM _G<9X>\MSW_7X[,%0 
@\&J0].P'E;O)/&68G<(92!@# H/2R12J_A2H@QB N;( 
@+XQIG?;HOI**@P*#=,E$+W]4WGVA)Y?;(M!TG.AJ;E  
@] D6PL!P37K9/.>*A4KC <^? ??9NHEXHO97<*!0$"8 
@1_K)]-M77IWO?X&!E'\T>C$*P\6K=#;JF!BLYW4PT$P 
@3N__A[6,B9LWA[16^BD*$B*,/]=7N9+'$[Q)<;..4[( 
@"!$?8F)1Z76G*MR7P"CJSO;A#W$ ]I5PF^8*K$TX'HX 
@PQX/7)L???$E.>JMZ([DP"JG" *(9N;[04U 0"X<K>< 
@;&EPAZC.FA ='36B:JG)_M6'S9#Y+(3?=":BP8#0LGL 
@L*)XG;6$;Z- LNK0I.LZ/Y3A[.!TFW#"=6'1B=56LJ( 
@7^02XE.HN)<J>+[BO<_W>/#T-3A"HE*H=Z]/!80W QX 
@:'^#DC_Z4Z)-Z$'[G!.RR6#)/NX1IC,#9=F!SF*O)GD 
@;+"PN5M!U"E %.&I29E"YU9Z_BD L5V CW<2>3]K/>( 
@6B-S_,T%E,B*5^-M4-/8?@O#NJ ]VIFILESI!;E7M5D 
@'MS]:M$68'UZV5I+ L?B$EJ<]-4EF8R/\W2_ ?70(X< 
@#O^UECD(Z1>2[ 6,:+C?BEL069S;088 OD>I&9\=@O4 
@]JH0RP*R=W+(JJ,#%C7,)DMT""EVSI@BI??IEQ0UXAH 
@F[A-9/]!POE26C"3'/WV9%1KXO= ,>+U7@HR>!"]M70 
@U,^<)Q%<TO#M;D'U@>K;;])L5Q8")(1(>3># CXA [4 
@UA%%@4^&%AEO3SY!1LX%K%< /]MU=@8_'!#LST \HI8 
@&DW1X:A)J5:A3RVEC3R8Q!*( Q1<XLIX[Y2(>?= AD, 
@YD<DT/7C\39CND+.-J?*I^9*RV^2\T$^UD'NHA/-YPP 
@E'167BK%4NQLWZS5NH%EBY^Z?^GSQ4:,OVTKY;%V*]8 
@\X%*T"UR/#R?LZ'DW3P<$?GTQ4J6LKP%RZWWV85? /< 
@DT<F&+.ZY)2])@NAX-?N\>O\/F<JF2G^J]I;2S0+AY0 
@*@H?:-]I_2,G=7=D@;YE1;"=L&%I&=;7<SN>.)5X>+D 
@'3V//N \]%_G_I]"8:A E96VC?_7&U5IA;^,MQWZ_NH 
@5;H!Z'-QA1M(Z""3/X$7MRJ:A$E[:09*J\(2;(]ZX8\ 
@?QTU6XD'%YZ00(0?<:%JO72_6*O5S3\]Z7(NIURYS=( 
@GH#I:D=F:(9H!&O.LD3"(,7^R]H+5J9WNI+6'NY\F,@ 
@TA8E@/&$=0UO,O_^0;QVZT+_790-..'B1+0DF.:;4M$ 
@3_SN@E.?HHFQB,>+4O+)*M1]M^SB*(7O-. =;#D"*%\ 
@]^K[&9?P_>4=K%)4'CX)5Z]C$F,P2:W*"L#67O4E_8T 
@MY@3%>O?<L]+^>8^]^U/4[L_.#2TX$;V#.C#[RI3]_4 
@Z(,?D^:^R*D6.V[NAH[&V/].%6W'/NL9RO9.U,+&904 
@,!CB)#[=?V#GI3)'<-+H,Q4,J/CZUF#CF,X/'R56<UL 
@K6IHZ78[#IOLB7DM2]"RG/,@Q^7>6D [:Z?S-1B5XY@ 
@RH"Z Y3_WI[8BTKYM&E9W/@^1PO7Z^)OX@0URFQ85=@ 
@%[UO>?8'D]RL,B&>>^?)]*!U(C"G(1'JCB/FV*87ZXD 
@DSB8F,<>.LX.ET]0"(!<.^>Q-9:9^#1#4+"Y%=J6;E@ 
@]_&3-RS:_P:!@2%S13V7Q'*-Q+.6+T4.G6"RGO/%4U@ 
@?)8C<O1MYF+P*=F!\3X<J;DO=@8-((VX\I_R8JHE<CX 
@?-4>6$*];WF%Q0Q,\$TQ,K>GV746;S^1.,E)89K\L^\ 
@\+3@NF*,V^6C)L?;!  B$-@ 7^J"+JE]YP.\E@ E4T8 
@,GK B%9_SU])45J)PX6J@L 8!'4OO%'FV@5(.*S'@*0 
@#-F@5$>]Q3%<"B&0=O8)>"T85Q1!4(P?(;&ZH&6**G0 
@PEBT<ACTPZHB=L,ZT./7]PLLT[,1A3K.G-:-<R0H>)< 
@DE*B'IA,#)W0Y59GM9:HUX]ZX"(L*'3"-IE,BJ)C15X 
@S-]/KZ*T$?>E@AN%,?)+H1W<(,$!:8@C8S(!N0XM\JH 
@)\8H!CLHW''[L=;E)F4P:UCT-E&Z[Z2BXCR_112XE9D 
@T4=&^4\2);*D1T"/G#2<,/(S5]:'X?;UNN/K'(M7%\P 
@R0E&\S4(1\V[_*6B/PB;D..]48)"L<IL43M&Z6ZMJ1D 
@-2*,[PN2B!<8=J1]T!2^X<Y7)[;<N9O_PQ18@<B11QX 
@,1'H!N8RH?T&]Q&GK(8Y]"LZBZ%&TS#QZ>0\:7IGO#P 
@LBF*M_T5.#M=B)#'U-R+B"Y01M+G?N?[R'-#D4A@@8$ 
@803U!R3.=;. 5)$7(>0I9T28V)J2#/1/=;N\#VB@.[  
@B#G66.0S_K #4?%!P3 1'O/__&#4FKW-4 O)B>BD,\$ 
@E25/$R<!+9VCHA5$/ _4:;B)&2,/P$YWRRS:V)CAG2@ 
@H*!\X:+IJ,BJT1,ZH1MD_Q>(JX88ORPM^AKXX@\<:M@ 
@R!BIK<S.T"8RA'J/LE+'G,FY\@NJ;T;B>KG37'))^Q@ 
@X#4AXD%U>!]>S,N(:7)6.(>GSN'\A*QS^7$7U[% XGH 
@$L.M6SJ0EVP5/HA/'(J:MT?C(;#6Y.AK:_N@K(Z"N(D 
@MU@^HV[XYBF63OJ@#)"37#Q?A;%?=4U[]T;8M#$6 $L 
@W6M2#) C/B0#:1GP">4WSQ1C6M@79XHHDBX!2P0D!7( 
@<?2,BX>^'E#35_'\06XY'*=%5YQ@OXQC\6J\!SO8]L@ 
@XS'N2U\N$)+\7(.)SMC;Y:V0@U39=SFW>D =,68DP0L 
@9C=H4##T39BG3_@ZV7&@#E\9\"CT+R"I\88HJKU@^/, 
@3B'P8Y"GEE-S=5B<!1C\!/?QI<B8APZAYH:D"=@[3-X 
@.'B\Y,-;]6/2Y?:5*FEBP.R:AEC2.M8.;XE06&@A&_D 
@@Z);M]YRPI( EU#P [FN4,87*=OP'+0_7@C >^WHX6L 
@Z/95" + S;+)PO.J#X0G8-K1U(BZP<?S$FOQ\D40HDL 
@A>>6:42\W-;&4;J18@.S0*X:/F238HC(,;RJQ(0L" 0 
@BN]'Q!?-"1X3O.%XP8-^A3!)@%QE1?QJ.$I=(0@7?(L 
@_W_<20MWTQ*YGMWU_[)8-UT[M^Z>=/Q<+)/H\I?B3:$ 
@= J;Q*S:RK\!Y8\<%K6H,9^O=-<T!694=F^,;#J]?8  
@TR&7LVR$=TQ^XT]2\#Z:0*+7=?>?4E!456&@ALB-NG( 
@Y+M!!@DFEP=MCT0,G:*UL=<$DU2-MW.C#F=#86/$Y)0 
@2=1CX"98ERLHOQGIR,_ZO/TI(;\0=G:W1C)>(Y-?*MH 
@53^(>2ZOA(5U71;Q -X:!*-]0;Q:%LZ2_,\C>P3BT7@ 
@]- =K:[7Q-Y&XL2E6Q%-P.(L'DR@HM5D0,- ]?-G,R8 
@[6F*3[@)<'2O_F!S0V$=*1A/.K(SDQ4A3NCJW6GD[]@ 
@4%.O%7DYU-(_7HH6Z64T0!88D$M=)K@<(>Y"D3$'PN\ 
@F>^P7FRLNU8$]UL%4SK\ITYFMQZYD2%.X=-5+W[U[*( 
@5N?NE[ %D.A2<<[R(:=SE# [ZH4H44J,T/EI'1$4Y\P 
@0K10AOS FP5;5]T(]')V^/A@MJ_H+J*1Q,UO3%;TE D 
@"279&V3NMP$!WZ9Q!]F2XV1CID VD,%^$&!8A]\MFH@ 
@1>7(%PA5YDE,842?%N\F3I.3>7/'XRN4%V'0:286SX8 
@%S#(AP4"<A/UQ 0".#.A/A-WS?='"NJ7HME:F%@$FSL 
@W5"";EDODWP6XVD:LI[LZ"#T2Z_PW(_8,16Y=4%VH@( 
@R?&X^:/B P#-/%IOBUEESHK-#B.)H-UY(ODY :+S'-D 
@67?H"Q@52G:^7'<EL\I9Y^(L_\IW\ X[M\L^RR<4V3  
@@L9('C1"7N WO(/N$\!?"_(,E2MZ #((_Q5P 4H5Q!< 
@=%=E(LS8Z<O=Q3A98\MW1!)S="FD2\( @I@LZR[F.SH 
@ER7\5V 0(S-83%;;D*(.X--2I)GDO*AD%6R;_FH]F7$ 
@Y4A*J2H1'UFG^-Y^[Z% HM&'4X*.!N%&VH)E&$NA+QP 
@),UUV52>E[HM7>,K%'LA7_3;3R9FKETU(52<'B ].Z8 
@*S_VUM))]A=:Q12(5OO^?@#2(2=R#J]UX1TX$S19G'P 
@,X%I#%2576>478$N4 Z"D=(2.2F"4O)_ VDR8V;WFSH 
@.]#5'J_YF:++C/BNTH7@BUIV#OU2#0%>2BX1:?SO!&@ 
@:O^Z93 F7Y]6O.CMO=3-M_T42;\J/$_UK$2?(9U]S'4 
@<) -MCKE.P?IJ8O]*2*^G@R4_?],+!?T%]GYN=%.TDP 
@\S3\G,(W3=^%'W7Y1IRML1>U0>.*FDJ(,X0R^!RV>;$ 
@PX<>/WW' :IWQR8-<%%[P"Y=I:K49#L2C_9?<R@\")( 
@NP.[29_> F)9U%(KB-C:"WTWH><D_. ]H_"\IL2!&MD 
@^ZJT<IC!9NPX]].R 16Z&0UCP*8X)-2M9B+%*&91OI  
@W#%$AZD#%>68+JMR$H_91T_1<2 WOA5]S:WY[Z"EP0T 
@VYN]QB[C6O/3@"(L1^::AO]<@]NU?RNHY#@RI[6>%)8 
@D9J23_2J-T'D%O!'%([[>B=VX=O*^\'VH1**:-,H]/D 
@*_X]B#@TEZFS0K0"9PW>D+D@CZE((-!025_T^49^=*0 
@9+4E\A;Y70%Z%H4'$V, .X, DS:U51-[Q'@*8('Q(QT 
@S0G:_K/Y+RI)YGH+BDM23RTQLZ%2S,>6PNQ,>ZO[?-4 
@4:B,Y^"E@[V?KDUQCPUR(QI=^3=FDP7:D2U=AVM=-B< 
@K$]0.V@Q+5,!MEBO>SEG:U+N7;GH.-QQO>N6C)S1Y"4 
@US#9Y#_%:SSUWS-*>(0A8U$$F#V0.2FFY_KLKT]JT:L 
@=MHP%0CBT/: HE(?A^;.9LH_*3HD.75$K'L7PS5-Y]H 
@+B5]H=7W7"21I$[!CL@I_W&MMG6_ZGCO:O+;>!BC9Y  
@>T\-BQ4;O1T%IQ>5P2[9./N&:D@NY/T1Q)((&E;D>QT 
@VI+ZTTG=$OLQ\Y.W.6"7SU>XG':-*O(6![6TDDHSB>P 
@UXIK0&T5ODT#"9230EBL;B<,ZRY"]%4S;87EW[/+K.P 
@XY0.0>[VXA"0Q^^I@*SC%1HS@IM)9.!&18X;K-H;^/< 
@N]P/\D];LC:_:*#\@G\+=!Q ;),HF1]E %N6),#RV;8 
@8>./I41_<6&WQHGA;NQG"IY:\G_:L88_RPF16&5@G_\ 
@K2BX%WUKEYYOZ7)SMI% _0BI?T$V5\1<<1>4RMKV]QD 
@_)@P'Q8XWR/5R)'2,$KSP 9"!!,6?>UD8G(55:KPF?  
@?&EPL?ET= BSV$2GH=3'40;QJ!!DAE5T$S9-:IB.%8X 
@M4KMLI>L+JPZP]V$@!:2_.4S^#T1/_<AS8/"D*E!\N( 
@4_BV$]'"[\L ^%Y%QVM4P+1T$5BU'[JK+JG8T#"M(F  
@[#1F<XL]?>VD:H"XOJF7JO5BI\D=CB5/D3+:$0\IEQ8 
@V8%YT44 )I-W3)BS<]/*R76<[625F"FPX*0QXI4@J2X 
@!&LFCYIXS31:2:1%,V'ADG R/D%2(FDMDUE-/$_T1"T 
@<=$+6@M#J'FB%R$"P1BICE,A7M(M0AU-CS:0FC&2H3P 
@J>6:]FLM6P0=XP"S;WSM.6$(X)#YJH-$>3$)$= C1L8 
@A,XD;%-Q;\A(MM&>7;ITW(11JL[%Y"UF3[HNTRQX ^\ 
@WFW4TY/2PYCU'58._2GK+'\,\;5FMCXFWTC:,/B",YL 
@8TLIE1Z%YIET0D);H%<,#;2G7\_/9UXR*I0=L5P\0JD 
@/W?,O6#?KX?27QWAIX=$)-".)0-\L<,A^72+)DE+B'0 
@RR;&V@;O$CMM+]HK;/UM]Y/Y#Q";8DTS*]I>Q!%O@44 
@6]D5UJR9*F,TUXH;7Y.1A)G;',^-X9QMW6(JC02Y1%$ 
@K:\2AU^-,U]'?>^P O0R1<ZIUG_1>);U96R:*0+191T 
@> M0"K(P.>G;3(<P>/F] $? D=MJ4 T[GKLSI]$&R$( 
@'M):T[TC3;6*F[&2?%YV#KQUU"SY2GJ 61'NV11"B88 
@7"S "$9%,SIT^J@ /WT L[*%S:]GIRO)(F\,6\5 1K8 
@\(6-[($5DQ\BAPZDFN ;^0(1%]@,8Q.V]SK4=Y5^H/  
@F(-9L/[>ZOA'[2BW ,;0VRS>!)' H8WS?&2)4?1N2\< 
@_=YY'LW-%VAV(^OY'>P+WTO4,93AF)%:L%=PC\L(S?, 
@5,1SN.<?Y']Q;_(P2STI:>@N@GIH=>Q0'<_9*60Z='< 
@<4H$V?PO7$UA5^Y"GL5A\SV,0\T[W[I"8.D+NYR?4E8 
@S^.>\.F8V*3TZO]RJ<1S"?]/[]XAVH#(!03LJS@L<5D 
@LU"VZ@@?>*!"C<L+*1/0KR.F;D_G_T=.,R)PIGC]E48 
@*;HS-1EEU:](482&A9.V/\//G711I"2&AFJIU@B.E!\ 
@NX$J*=Y;*Y!U@=PM]=B^X&Y>T<=#5O# '?('^0F8Y)L 
@?W/WA8B%=,$/1]5UU5"S9=+9.-MQHCC\Y*T<1A+LN5$ 
@J>95G6C(L!(L-E\G<R*.Y"(;)M,A3NODDD8BR<7T1@H 
@.RNTH\=NGS[$]5W+!+NZS4?IQAR)8,Q1?'GNY!H]\-X 
@MU3MH(]ZW1WY!MU_- T^7U#$C<^?AE9[Y1X;86<S1VX 
@6+,4)O;D'4UHQ'1T(CLO_DING(NTP'UCMZ4>XK#6T#T 
@VQ2%^_;7?I-X,4,EZIBJP/S2!3%K0K1IKJU:CGG^IJH 
@A\1XT$U#-O2$FF^9LU#K/8'E@T47JR#2LM#,4V8>;WX 
@V,%'A &A3-48^L%>GFZIH].KQ%/$P2+E,0F(W9N.:T$ 
@"*TVES*--$,:LGC8:+4](AO!C?<^&Z[9"VSZ)[5]&/L 
@A9)EGJ71DH!9[,W=JL3-QLARBJ>_SL=&M//%-285UWH 
@!R+&PE5B;:<K!@I!&\-_1U?AZ^3++N:RA,7LK#^GLCX 
@=J:%"<;3J9"S)S.0OR7BL1'W0W69T3;6-[N/YM+4])$ 
@\"9(>VDZHGSC:/1FI^?Q-MMJ2(K)0\\2N(N?UWQ@56D 
@#].?#M>4H5#*GL*$>Z-  (3W=CXHK$<-#4X>$O;W.T< 
@'J7LP!L1G8?8.43V?A7O<3Z.$"Q#66<G-'S"[SA8;IL 
@'6>:S6 5P';A6DW!8, JAK7$".'I> .BKL(U*WPE*T$ 
@ Z^]->M5UG.T.F\#3[0AJQ$IRAX IV>=]!MA^T[L'0\ 
@$R#^9HA0<YR.67YNK^ZO5T+O3OL\*)V&&O.B.US:CU$ 
@RHK^T\HNALR><P&84GX1Z,F?%= 8@+O'N)4-?]O_YY, 
@>>X3.J),TCC<C*)BA>5.0\G/,JD7N50["NGXIG>.E!$ 
@2\ADRO ] 4; ?UD+<'1T5N-316_+&PL6F@09V#Y">+$ 
@",C2I9[/3GG?-P4*9+X92&&<_\YZJ*]2,?SH#+:A9*@ 
@QDTCAK!<#@F;RL^?_A1! 6/QG>PP(84I)4 SNH5_O&\ 
@NW^TG&1+&/O*. M..0E4%Z00#M=47\>";4RBN\B?60  
@>L9)<K)FU4NGK4.^!M3=Y02'P-,7U=_>&UVF8EES3UP 
@V)PN-YIY)%U) H\S-PTQ)J%_9Y+7V@>K6O\VYR8:]LL 
@O3#1$@O*V98B96[WB71M,G+^.Y*U;A5^SD+JIG)MB<0 
@]YCPH(;+S#IW<O&XL'\ 9C@U89>YTK(<TID:4@]EU=< 
@63\%S@60[P)!JFBI7[C/@DSF+S9A7N,S0G),=I"_6/P 
@]T?10^CA:]FK*VH)K%XN]WJ8J:!6BI.&(![^_0:D-]$ 
@%0\:.+^#(S^E<NMHFH"$,6K[+-2!-_1$+#9XPAH*MT$ 
@?=<(/W/6[YMMAH:;A@,+/,#=W[^YH0<Y6M$Y1#M).=< 
@&/)FE3%K;,J\O4RR.==Y<ELM33'T0.$/Y&_"X0IKHX( 
@KAS9".0:NX[TB)MSYR _^:L?%Y]5-M%=8K=PUHI+8QH 
@=OPZRM!MVN^Z]P 5L.?'FUB]Y3GRJ0CW^K\ 90?X18@ 
@A=OB+N#&?3F2P_1)N.OXSW8ZDF)RP5Q)O1K,9=E(M2P 
@K/7\6GD3S$KC6-I::?+TY@RJL_^P*NY]1!,6\PL -K\ 
@U$]?P*?Z%D^EO,?)G57UTJGH3B7;IY*-$Z\BF]M'\&8 
@2CGI1PG09OTLO[-"<'LWEN.K3-@EG_3.@B0_TF$CM(, 
@FPR![QNZ)<(EL8' R%*4,9@%N)_5@7J%:T$%.,CL]"D 
@]&#E+F"#/;O /6-QX^[,FJQH:'O"I:NY:@(RUYC077T 
@*L?T34BPV\\"A7[YN_['8O2K$!$*?@FQ+UMCWQY8[#@ 
@ACM1I$5R71>.6-E-*DR?SZ^2>2]9QIC9W4_'M.UL>>L 
@=6UTX&ZX(N&8;0\,BF!3R^C#L&;/IF(XFAV JV8UTLP 
@?L ;4L&FF '\IZIHE/=D2;2'W7-.,53K(O'B)Z]6%XD 
@!]PR'-\:6^%Q1(FA?.FV77'&[A%5%]@N1[AB1:D)QT$ 
@\)C+ .;'QP7B[H1KF_^BNB</*^B0GP41C2]D)MS .ZT 
@P& \^.0%#!L_@@)Y%W<F(KL9KK<\),V62H<FC 0F'ML 
@;")6\+ S.ZEXP.XND\3W0VP\7&[]5#$@[)ART9VK&J\ 
@>IS=I%T-%4-$_Q0NP9%8HBQM(JO25QO-:3Q;HAQ9+F4 
@&T+$4U=#O:RC#&J-EUG8#_T9;[3M6S]M*)5TE!H_@#H 
@OC':(),>$W^A7(+6M/3B3C40_H-%IL<@6RC.=5%?5$\ 
@!Z79CG[V\&<&1O>S^<D(2&G6"QN7!7WG7+ UFHBFO,  
@\8F<<?F&XG%>);WN#NC7* (WN*NUZTG[0@V3XS9.(-8 
@WE6U&8\Q^D.).X6SMPKV,+BX\G94Z*=1N+UZNU@HFYT 
@%V+X@M\+5/>J5ZSN.T2T+^^A/6 %6&9?.H$A$<VN%O< 
@(796]8)[55146JTSVJ<<Q?3"CM,S.$]$^B.N_#0A(-4 
@IYD#0A48L!\6<"VE*,PH(,K_HOD@* /2I@Q]5C:A'6( 
@DJF82^ONG#KDQ*C^J@UF*L5)(H5BSCX;1><)0>8[_&4 
@4XZDRIB3).T(=:N1EJEA7R4Q RPG7;EQ2B53#I"Q2*, 
@L')#T;W?Z"QX&?EG7I3IWPQUL/,M]G:P -K=WP21O"( 
@TUPUM0T*.ZLPQN27^6S<*,TC+&\$R9L3?\2_&TTBZ6D 
@3N008##$B%1V$/#% :4, UU% ,L QH>#K5?<^\E> 3T 
@B9-0/:O>1-_"$8U1/'H4A]A]A-5R%#7W1)#B,4_BZ'@ 
@OV696;KEX[W_(D^C/4F.+#M5Y35HJQ8T$0K6X[(.:/< 
@%DH3OIQ3F;=VD7;97#@:(=CB>'T;#P=*T."8=;:)/3X 
@DTEX>K]&]H#>3#JM8A>E'S;ZQ]V@><84#!5DKM=STM< 
@DF-E!QF((1$B!NZA-@J8L5Y.C*H-\LJ+Q]'BMYB&D4X 
@BM0BMB@2;HC1V5V DM+SG27$NULT<3%V=HG[LLYPF9\ 
@*L@;*?78\UG[[S) H=@"7%NM+]W0"%]8<[N6V%9BY#0 
@PEY<YS(-E"J$Z8?]_]"3I9 R!=0/EJS/^FY,_@=VMQP 
@#V\$>M'%YQ/R2A2_@Q/N/TT0,:7;N:H]H6],ZV._#3\ 
@SN4J Q^(,C<C!-\8'6KN8^D6(>+=A('&[H:O""/M@_L 
@0EY1VZI^1M!:J$>LJ)$V5%Q[)-BG;!E.0F7,62<^U]( 
@E$I^"YJ$F78X*T-J,,+!,<6XFS^?_+>8E93HALDOGH< 
@"2^+,./NF;^E(FD;P.;52CSTS\_%3;'*4O(MGAL$8:X 
@NGPLGU25H?=$U-UP.4@&R@J_@/BRKIIL) ](T"E69>, 
@TB:>"?DUN@3$I<D7\T-K]&N&G$MY:1<%@6$RJ1+-W*8 
@<<%3ULY*F9DNX)[]ABIUY]N/Y[QT-H0]=9N=1(BWLOD 
@"A#6STBI3:GTSCH\,NCWM-2%<9.< :4-.S[=[)*2]R$ 
@K6X:X;!_!VTW"GN3],T1(T"%#BDN:FIJ '&8U%1V2TX 
@12%W;DBG3+[\(97_N@W!I'1(MJZ)'=C'%<1 JG6VW@0 
@S" NU[:BX>Z[S*<7^3L_.F67@Y>LA%,ZJ5Q"[7.$$LH 
@/?<+^:$'TOM#TD=*U9H%$2WM5+&C%3M(-0:9V0/$M , 
@IROR^T!5+4K)SV'B<1E,GJ:%H,5?&C4>Q(*/Z$1!#0\ 
@"KU2P<:[W\W0)=E!:%-R^GVH(?^;("<R>_LD/NJ_K"( 
@B!<S!R)%XHJ J$1\HI-+P5,M!$QD?7;:WV-]BBP[\48 
@0>PWA:-JPP\@55VQ9O\GE,IS4W97@Q [HW6'IH/S@I@ 
@=,)!Q<*(!Q@(W?+=!RM-_/WT@^M795SSRA498I''U0\ 
@Q760I/P:==7@O]I0$@C++0XDY1' RPFG;S!9^0\:Y/  
@X5=R[$S==.B:OT/=M"Z>AZ-3J:5@:2^UANJ4HE!(BFH 
@;%#F/ /<&T5/NQK&3CR3#@'KW2FHW>1Y5[J&S><50IX 
@R[Y4&U2D!;,!YRW!&P+27T..RRW*'EY#33X=@M48/IP 
@ >1,G1S9*3\7A7&_W#;==K+X:]:LMC,I^IX3#KT>ZNP 
@WKM*$,W4GP4IQOF<ZGQ=?%D2=!<?SX[F&K7$6,J/Y-, 
@@CS5[M;E8L'(##6TFEHEHB6.K#I .U_#HH@;JX5UE]D 
@)]@0'X6:*NV &!1POU^R0K"Y5-*\UWK?PU T,T-4\XH 
@6^Z&:%-<O7GVNY5NIZ;P8L<=PM@>VU)J5S[3_/ZKJT0 
@!5M"-:@TL%-S:5N^MG>E9@+SU@RNB@$@C9-1]U7^&38 
@D@G_3S_8J?2J?IE<#TJSDOO?*QTO#Z? GH6\&:E1:5P 
@5R]/,$%=+)9OARN2M'PN&;?K>.U1*I\;D$7GIUF8LKT 
@Q344='/%QM^EE9J#H"4[\;M>45LA7@8@4!]:.TZ)F*D 
@]8JXP<7;GI&-5CANNNK!XK:V2M>+@#32(A/S.B!C/5H 
@$C!)\PLO#PZ-8.MX3M(31ZNZ/J_^>1=(5VH;N*"9F.H 
@"S5-"\A;VMP;U[^;QYH\ML(]R0=.2G!EW7\(N\ -'TT 
@X-S7>@UDT^N_/;XG,FU#3"!3\UQ]!U5#?W]?U<TURG( 
@EEC.;KH&>ETB4T/J7YNE[C:#HAHB;T."<+7H:[H]\5D 
@ !^J]\E&GG P//=N\9!'VWW SJ0G!>*.MKL*!U$O,44 
@Z>I-'-%5FS92M@^JH_9+H$4LDF'"K7$3^H(\6T%1;I$ 
@Q8S7%B+K%H9BM6YHO9&YF1QK" /KHD6U,7SDJ8DPNP4 
@WF]%#_A/J ]MB3E8KGZPQ]$M:L[/]'[FO"=RNV-P*(\ 
@K0T7!@<3,\G7Q7/WQ= 2G#IX5)B,#0/$%<@--$-/N;L 
@Z(7:<V=.3 C(YZ%CI;/##ZY@MKV@L<8@QJ-D- -EE0, 
@*RN=(X'J83/4<N(5D FRU^E[)48\6_-C<=\T^!/ 3_0 
@VBHNR>E%)0V<)!G_O^$L>2>]R^/:P^.X!+,_PXHX4&@ 
@B,^ &7^;^_(^DH=M7"A3:B/^+"&$X91:JLZ:7I!F;#D 
@2(;$I%:04-O+/%X41\&R1 ABGITW67S:-N,")/P& 7( 
@;];X,.CKXAJYB,HG^48FZX7BB8"C37H!,]VY<5+3SVP 
@?3P1'@:Q(ZLI)ZZ\*PW<$&PVA1M^=TL0DLVP)HF/-[< 
@-<HL:37@#7R!Z"3V.NYM/WC:/?=Y38C#Q6# !D:#G:T 
@J/)8TCO6AN(GUOKP$>/M?6\'H76R1?GWACC/?D_^;Y( 
@,U(SZ"RK9-[,"F?A3Z0FNB-)F=N%0M/G("A[&:FIVJ< 
@[Q8/3293]XF4M[M5Q$ TSI,+"S6>>I60=.E\_&-!QA4 
@^/I,RY]Q>GH3&Q'>T]R\;E8]VVS#Y%LO@=.%^']GF.0 
@D$T+LO<43G)-+##7J?^ Q@+2I1U3KW1O>7-90%"7V4T 
@./GBN"I1]Q".1_6MSY,=1L]H'# _EUK6[#I_0W%7/+( 
@IWNO@QEH6'0/_;?T/AY0J+[9J"WA=EGG.E5XDZF'/1  
@*;#<X/L0?7U'J<6'Q$MXQR888/E9O:*C-2=Y"8?QE=, 
@:;UP9#$W6)I"%&O;S.TX&*F7[8:QQXRFR8E;0M;%5_X 
@4";6>*3>(\?.KT>M"\AL1@WE@!_ -G>K8S_Q,/8CV"P 
@+K#C6(L<;@+L@4/3 H@_48$7W-Y?52+6@] _%]CG0ZP 
@]D7O]+@G5?4'4!58.[BN?E,Y]C^+-Q<MWMLA*/6#>!L 
@!M8[L>$NEHC*;UA3#K705">$#"M *SQ]>F:<\(+R_SH 
@;6P07W,+L'JZ<6A""Y1:4(*#Y$<G!]#!^:54\SM#N40 
@32;T17)R&@WT&:S=4WY3UYZ@Z-^1I^/<&(--V 7HL+< 
@,FZUA;*U%G/*6=T6<")"-<V<3>(]D.(GSJGYLO"HHD@ 
@JO)9M\ZF=)OXP@]N7!2'*=4:GS;VK9);FYPX60E@[I\ 
@I$2@9:E@UY<\0<PLBQP=NDS4/&5!IA=@OCS2#"XM&:4 
@=FK+N-@\\4%MK>)68[-"VC[  >8?NOSX5<P;>O1/(08 
@:9(>DG8>QGRT#<A]FQ,*/<-V)$[",J#"*-WSVPA$54( 
@2!:4=/'NEFQRV:IUO+@?R8SD: &^&[0?X"1+* @$F5T 
@->2<;P1"H.Z5KC'=&)93W)TZ60OW[!K].BZH<;%L1(4 
@&HCQXAJZ=&-\ J+=B/M(?&C*PG752;GZ"&C+Y?521K( 
@6U^9-<H0@JT PBVL(4,+)>N&#),- BK<S%PL(\_JST( 
@#8/$WE\<"?LS,L>[S?3MZ6.Q5+9:K)=@\G7/8.?32N8 
@]8Q2]^81;3@P7S[:+4&YS*6%HOW3>,@4:UDP$C@KQ_$ 
@$@(EJ/*>Z34B89::_P&F*Y"M@9O7V3\$06?<]AC'&HX 
@F^/WW0A!8*+'#N.D!@4_[.7,63K3)7VMERJ0LR5N4*P 
@A>#U_+!>2!>*WERLD14$V,8(W)<UVG8B%K=R*6T=;9( 
@ZPK#_:)MJ.84(^'Y(X#5FJ!Q_1'I+5 C@WOL,PG,YH, 
@M.?,\_T7Q*ISZ,B/<&PH/.ISU%<NQ_><2F[/%_(,!=8 
@&N^&LO^7ZG;U-89#K5 L!B9X$BEQQD9.[UMU(^S'+U8 
@CF7:#2M(T7-.!9Q%M[KRUQSV+$F#-R3/JY^H]%I9Z@H 
@YM!*(]4GDP=[3!V]N^8>9Y W%T1:_\%D4;UY#J Z:&X 
@ EIYP1D1@(R[!8"#?Z.VA4S8)UB^O_^I));_G7.SZ]4 
@1!.1\_MVD9_,9=3D1.D#_E?*PNPKGQL$>W-!6-[XI>$ 
@'N R(6:=O[6V_>N/%OIER%ZN37[ZMSVPND9F,9MJ8*8 
@6Y9T3Q$A:Y2#HV671(G)^I^' D+>0C>CZ@D1,:W;-Y0 
@=,^YDI..9LB2-M&*2KGZ0!V%SA(VT_L:4"!ZSBP9#=T 
@98VK7,VKX5^.I?*S=;A[1^+;AQU';T-M"!H,"+OO:ND 
@^<1KN#VA%$D'-CWTS^/M"PM'XER-5 [,2?3'_3$PE4H 
@L2"$BFMY!?&W'L?/DM1*#VO-Z'A [I194(M)'$GC(&8 
@',%A$SC[A\]I[C#O^&4C3S0].C_V6S7J=@"GCZ:ZDQ, 
@RX#3"Y2P5ZV.R7%VSCG\>"G36DRHB[@7&TB<$DYQ*'8 
@.C6D2H.X6AHK$GO)*&$W0T$^US6;AX>9)_T<?6VERD4 
@0H5(?,P?T[V7\9'/[+R "BZB+M 7MB8+DX!%$[)Z)U4 
@2Z)MXX,(U&NQ5 LRE']#F*,H(DY^\[-;=*GQZRE01TH 
@^S2GC]*IX^FA'^,\E?WHQJ0/>(UWRG[W\VCMO2*#C$, 
@^Q3K(H/%T<;QKZKLAVJ6:<JGL3'N*1BNI-=OO'AC3T$ 
@?"O?,+KX5"#^4UOW+PDG>W&FX6!V-U2G)P2H:9 A,-0 
@?SP+A2>(M$'TB3R,A(E#HKLBNZQ6A"''14[]^8A>KB< 
@*ZHD"=/C$D;,W.CY3^>+%-CYE)C), K7MV[L7-?S>I8 
@$3;6E+\7=J(E+[VE6E"!95MVLSWQFD^H1AE02N^$&)( 
@<0(Y;*M5218R0(Z.,2DL[0-.;A[9;<J?0&BN@^S>4R0 
@BG(@.](=#6TU5*616*BHSWL9Z?:*> ^MSRW2)^ -O:4 
@X*9JXUZ+,\N",I\??<QM'K:!L:F^?X.-G%;9X*A%4/@ 
@P&"KF*1\\! 08-V6]MPXE3>80Y(_B:_4=?REF?6[&-4 
@4I^FGK)_@^2%-JI2%J9Z-AD5?%%$X711^!&(ID/,+6P 
@)F;A*Q!;R,+;D82RH1 KB0T:W?_R& .;9[Z=G!5Z32P 
@9=+W *SM@?>SI1?7B-,/AZJDC:X^8I#]+@KG-@V)+N8 
@".?\%@?WJAP@E[GI$]RAT:^M+S4=[;IM]VTH!OO4;Z4 
@ :3SJH=X4I<=2@5#OCRG!9Z38TI"MN<HNRA1M'LT?:@ 
@!&S8E*ZP)W)PC28I!Z&Z 0=<G3"OT<TWKBD_V=6SUUH 
@3RE6:W==E]Z>KVVC."Z:ER36/+3ON5\CY"Z[AB=@PV0 
@BB5<1O?PQ9QE[_D&[N;-[Y@,D_OZ!/R4NCWD>H?K3 ( 
@]TZ.PO5-57*UWI%Y(HE'9Y_4C(J_\NO0':J,QO^:YT$ 
@G5JQK>>%I;]]D3SFM;2<X/!_D;;W<E14&WCU*';+-VH 
@6"UH^[:LS>@$X-=9G@6;R9:^?R7'6=J92820T!D"5]  
@[Z2:MP6I>M5N8'34+N;R<*Y/OQ5YO,%U'#K0S"W5^7P 
@<PI1$')(QE^NS @?23X_=:Q<&CLJ$8>SE 9'KX#<%?D 
@INY&SND#B--LK..E0K%\!6/6YH?#YUAG<K?QI["DQ\\ 
@\HF<-]K%I-[0* <33"H=!S".4L?=3!$ 1$H'&[;+R0X 
@B2E^DA.(G54_*'UU#RZL"KGS!:@&'!Z2]>]97H*BC(D 
@O>J=0-C@&\*FWL(('MF258='TE%#8>%AP^;(:<?*[O0 
@R!D(F=D0%8'>J$"5Q]1:$&N\\VU>;MSHP(>&^F8&'O< 
@4K !"L.5U\^]\>L12]WH!(_8\0*#H\++7@\4^E'!P T 
@:)\T>,'6PN=':=3@R1\CE3+T^SKXT689^ER2@QNEELL 
@("00OPCC_^  ^,U,G=CQ;@U3%2O#ELA5CE+K/HWLGW8 
@B9+]7BIYF(@TX&'T8! ^*DIY]YJ"'MY]GI= \!.E'_X 
@) _="5QU$%2Z;EVX=7&1JGWN=+7+UYNC01?_:VV<C6$ 
@D@/Z/7U4]VA>D!8:V/+?*ZP"BPVVFRHYUS_@>/>(70L 
@#W<HU/A8P<\K.&!-T2CZ8$XK-?UANGYKS0;.*L:1?8< 
@EM:JI]"H*&8%V[Z';#TW8WKIPWT&K2.C532!X-R3GC\ 
@4,]^R>>R$*9[<9W<E,"1F&S5G<#]Z%X\6.I:S_V>PBL 
@,C7:W4!E;'&U;>OQFJ(1=J)0=E#N^!Z9+?54C+M. R4 
@-&;[T].M6+W+!0,"Y#"X-GY)DMZ,L)':R>F]?H7KLDX 
@\?>#_;$@9&[5JE,($NYS[QVW\4PY9FF'?E!GP)HR@GD 
@FC$DHOD-1) T&QQ>K<.CW?(RGRB2ST&.#(>[-V8O%!H 
@#49O) :"-U G_HWVM]\A6JY15/AN-/EEHJJUS-(5TIX 
@0!7JC(M2<-([/973+I&Q,L48\0ZRM.'9")K>WTF8ZZ4 
@TTX4(\OB3%C S"7Y18F B/$SW[)@/,\'^L.T@=F0$98 
@IH",<695^7\C_>,K:D P>K0DD8X<UF9^!SK.3*5G,9  
@@6**GJ"R)T@>37 \@_&VQK 8-E>.<(QSW:U+7-KJ[.$ 
@#':5G(TXZ<NGO,HIM?N1N" +B\J]14M_E5:QG0,JLG< 
@%%E9!.D_^CV+PL^:"%LF[:?8^7>U_ FE9CK!\(I.UST 
@M6/0W0WP'WW^6@4Q7B$YX54Y\=BU?GU M0?*;?&KW<L 
@6!/\)XU?5=S;RCHF)?K_'O@[8 [[#?4Q^@A/M9$TT<  
@4]%_],/O#9@YT1*G@DJ6/%'$#QE>]"T<S/R_1HVHR.P 
@FD4;+@@ED\K6]@5(G@5:-Y2:194_).L&>-M%Y_;R,"\ 
@U4]+F>E)<]APU1&YVT.@7W? V"J$*NLZYVQ'#=1[&., 
@G+WP>K7+P#S2L5=#K-H/G45E7+=ZE32HV?T^<^(=D.$ 
@& .1]6B3F&U"V\)G+)5K&PM]%YK+M,JN^-$!XW-^4I8 
@S54T^3:X46J(I:IDM8&^X$<^?)3=Q>/E"_T94S!AI>L 
@0+'>V$I,K&^6.>1"BPD-)*,X(IX8.R=GCG=,E1WK72$ 
@M+UF)\D2"N?E1=MYJT_&@0X<(JV8WJ1/-WAYU/&E=2  
@M+/KU>GWT7'F%2WL'X)#)]]SDUF2[60,0Q%!#X__U28 
@.V_W%[&'$;_^D!F+<.GL;\EC.D6<ZPQ=H\EU,N-59EP 
@#'HIRJM/J,NL&]="Q$OR9:DR,9=?Q(6H8;E0M!GT>PT 
@]-Q?40GAM/42V8<%Z*IAT13XX'(UB*JWD:/,*8B ?N\ 
@-_W)M6N>8X:1[07556AHVJ;=0"4Q,V2;LW.+<*UK]68 
@A5VE\CH3Q1L?I,=R*%"B0 5-?_D(3,&0S6'8P=+Z"S( 
@@U9&I#'[_H![2&+W44#ASW337[1C-ML'!B^K:CSD2'\ 
@JGY&MKF.P53>?WSPJ04MZVRY.($@Z.G8_@Q=T%O*9_\ 
@CR*<MM%.M0?&I!9J>!II,\*8YM<)LBM1W Z25;)T7&  
@."AE;OAW;(M3+'DLMTJ\1-)UAA.*Q5E5FP2W&"??YE( 
@X/-J)($SX7@8LMH"(H57N<G_H ]@CL],Y1T)C<6[&'  
@<]A&LF2(LT&>TTF335@X64&O'M<3M-[9?LT/W(:]U24 
@D8NR)SD>FNKR]&LA^0^BRC91@S6 &^S0N1@=6I?1&O\ 
@![>3E#BLK"X'\MHDUKPNG)J6E!6N'?X=NOK!O;O;G!T 
@G-(P+# :EI!5NA\@#=;;KO %GG<0&D4+I7OJEZ'1T&T 
@B7!0U4MZ'* G #3NHE;-Q ;&F9O!N<#Z#91)Z*!  +X 
@K)A*A 9Y$^^U=*('%#!))B&#\V\)?\$MSIS_YN?V?]T 
@[JB16*VD0Q5"G'Q[7J*_!Q_?Z'G)GD^7L&!,H%S$,44 
@4XO("U:3'/-1'A!P_*I@EJ3K.=^-R<2SC;% -[E.);L 
@6=6&?.><BR2LA'6]<Q%:<V!P#^^V!-P*D+!4!,/N._0 
@BU,0,M/(QUMQ*.W$(F',.%R"A+C68R8PS@"%7!/?)6L 
@/=OM/=LH< DFJ:\L$>NOJ**O/FW8L?PR+ 5.+WEF WH 
@0ETN-I0V?"R5(L^.<OU,*D/]CX)K&"NO>Y=:"MAR;6\ 
@$:J3$]:4 GY0)<\Z]\R"$*!Y8\E6^3<I_Q@S^^WT;%H 
@I_I+W&I,)?WKWXU?8.@_W GT_ EH?9,/.+^%M=[D158 
@?4Y'.^)T/,^P&VUX=9)<)S!4WDM+L^B52:3RP<\F 3  
@]J1Q'OB57#[LV2%T+T.'\Q?Z( 0Z/6G J05Y,<J# /D 
@.^'VMH,9]K F,J'CG?Z)@#'/#344#$2 8MRKRMD]M ( 
@VX3"NSFVZ>W7IV0E+XL,30WR7_?>9'F%;V3&1%K^1X4 
@_[C(SL3CD@SL?!O$U=BL(@ZE#UR5;?O0UDWW!^%*(7  
@]^WB&,A$PCR9HOWC)UI")_UP+NTX\KS2<OYLE\)!+T( 
@I-S1!0FIH*]4D"O-85Q^]!3%=7$RE!,I\RB\[_6Z<#8 
@VD[7@3BW,\ 5'3F$;;-5":[V,76D:)L$:5=HX1846N0 
@=2;8\_=YMM$ XOP)WDA3P?Z?/SR'0!"2/[<[YG3ILLX 
@T#/F(>F:A0DF&"$R\2!A;Y8*!.?:!LD96* 1RUOX.64 
@G?*^=1*]6M)QEB<:[59%!<]A"*6C=TFV.YKKM-]%?7< 
@(1(-ISM/&7YNCE&QTBY[K\N4E(S,%&&J!=!+B"=%P%( 
@XHK?@AC;QB02/B]HLT\,RA! 3MW@0HS8(9O#I7%:!SD 
@2KE!86%!D[@J5YM;;/#!TA(^ #M[59MH4K4""!*:P.T 
@^>!4#W.E B?"Z:Z-&_^G43*XEBI$%AC%9WP]6:BOV.P 
@9<7/R_V<P%K:[NW ?MCOOP)Z:)O2LVXPPW3,5!5A59L 
@GP23+U^#QPU\$,"31%#=<&REJ;O&;GYFQ8%>!BGG3LP 
@BH@"U,955WYWF&T+1:N&PH@!:7%/1XA8$9V#'87-CXX 
@=!!E&PZC8*?][%/.O]DY%(HUN=2%#MLW; &H,\2-W50 
@(V6[E(00@+Q;CFBS*34'J<^(D%D+/AEIYU8!S)ABU_0 
@F >;KSQ:1;]8'W<;#8-@50UJG,R3Q);=GT]XSM@]NK@ 
@R9F>E:D4OHS^A<\*JR#LYM:?.R)O8$@E^X6A-]99340 
@SWU"S_=KW@7DGJ/PT,MM0E0T>*D8++=G[L^2(CH\8TX 
@?B"D'QL$'_<1E'-4FAG(8?@C:_,])QE[KHW-9B=K^ZT 
@WIJ_ZJM6 %>0;MJHR:YKETZBX@<$H:(E&\M_)M]J6YD 
@$AQ_>NO)P?LPDQ!\$5#JE+Z?\069A6:GG#HMGN7T##  
@._O[(D3K]_!P/=PF&>%CQOV-$"Y@ T&S5/20$1++U\, 
@Q4/ZZ$!5QMMUAU,U&H^@H")FY+$I47K<)F2C:?1*55X 
@5-&I#)'@7Y"RK#R(94?^3U>8K,L5,"+ ,PI:>(8Z.LX 
@ST'7-/(D(?W@V6GJ>_H\[,W%HSN%MEVE20!4<&5'^/H 
@]YD+Z.(-*]EST.S5;9Y)+^7[A^>CL%)]$"PMMM0I^KD 
@OI\GE3Q%5N2Y?A)4-U]$AB(I11GIU\;M0IJ7=%T0C>@ 
@0?JB_FG;L/R3H'I.Y+>.I003R]2FIKR'E-2F!?TMRKL 
0WR-;N%J/(DE& 166!@8':@  
0!#YTW?!GH52Y>:OX'WA/-P  
`pragma protect end_protected
