// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
NFYbNUfkaObonSXwz19bqNeHpBPrQ4ng1A3edsQgdCf0da/5lWVvn5NNNEUii2qZjjvBc+wFMfXM
HwkQDKKTip0IuTRkMt4tgjTQmw4fBR3pN6QwrQRPK++XgmhtuwB8B3B9DErOsBMtS6zJhsXQ5f4v
dja8Njlq+CtY7dpbUv/Dkw0ySBPDzU4loO1uvBLvu9vnQw4GEmlfaRVbavr4l7f+hvvTcqU7z9Wc
nFnqFUR41tdZY/Rxsodxgk1AztQPcTl1gsqEf4TJA73DJaLkP5VJPswIaTUS/kF7X4mDX2ZrP69E
Xt2UwzOZZf4B9a4japkakHj4880B0zhO+56LbQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
6MEIqKTYeTiWFQ3WpVyVUn5/IKC8a9VPMlLGjmo47hU9SbBZu3VmePNgR+SHbRTMKQAfSFdM6TYg
tgKfe7t+3ZoX6lVCz0Lo2lVHa7k7OSFq0x8kM0CQ750gWs169ErcSRCU5rKqh83TcGLzglxhNcdH
2ZVZlUGje+jgz45Pbz8InKUrU9aCvVGX3hQXqj4tfnhcSC2n+u1nQt2EFglI6h5D6eSUHyJ5txYA
002UPZOMcZWuXqxZmKCLyA8wNXXkcM4a0VkYe2dNO8BR+di2UoAJ+YSH2lVrAXqlB1Hjx4oVc8NH
qA1766d2zCOE9QZfxeaM3BDgkYkPLp2h6QNeKxkjBzXE7eBgJg61ehAiSxptbR4e0GbyxQQFMo51
btWGasLos2Y4R+RlPa6b8Zxbyi09nbdTy3G6i5LXZGB0zONndbJ6BtQWO3fnnUCdfrvauvAN7cka
TR2alIUOW4QbJL5+JW7OiEuV95Ac7oYXIXHemb+wE+95VUIDk2Qxs92zhWXs2k1j3snSBHvVuCCa
PtsJQS9yn6+CXcnNiEZHZXTMnpmXJaI1XQ6pHY13MZHCzUJARQ3PDA0mFS07M70SuVXfNzEn137h
YOhNGmYYBl2le/Dv6l06VlDVvoO7HdK3NxBugg/4JGmQxSXLbTagaLcl38fiuFb4eQ7YmZ/HULww
q0sLXLHHMraebdfqsjWrr0ShFHCfZxnOdfEYx4pYhOvxkz6std0J4tOd60qSP+tAF39kIfPzyg0D
8ttzDBrYLzDE9NmY3HjS0tV3nsHlFwnUN1WSYBKb3MhOou3RlJbacEhCO/JUsyITsA3UM7CcilQ8
bePffOibYCTgOH5xIBHpPBlkvD9LFkms6+8bw1aTg0oOX84ulpwCoqXoC9KMYUCjrKwmxCZ/iDc4
VJ1Za72W7WBCnIaqaRd1O+bqbPniE9Zao1MvD6oWi19HMYh/lDaJR8/iF0pc4d9tDfQdlClP012+
PO83HVmu4nLO3nTMZBmfzCdaTfYPogEijoV3gLc3EtrbWcYGjgzqBdoxry0FbegzTekhOpBrMwTO
viwYXdq+fOSl+IPGyOdcjclF8HsDkoGtaHhBw4tZ83Rtdnfvo3nnk0x97czQyAZQpyIgKbDv9tqe
GMF62ezl/jfgoIKqbhVFt947FzQy0vDdIStLCJ8fSbOjGGmkqD1EhJh31YB4z7S16h3P14RvXDfn
rrGXWgR3PZs3U0TOLTbNRyXspPT/MNO9yrNh2IysgE/b0vnJOyMkgqO1BbIerxqEtKskHmEn9lKU
vRamlJyRYaBcSuuwZ39BNjSY789jUWO5idKtSVt6fIhlCblHSq569cMwQZDLwA46kfH7xyRD9DnN
NyHWgjfkGUhF64Fn0XknTm0nJIzqNkq1xKoJlwH/fYRxIUkUctXQcbi4h0xP7cbl/Zw+zqcMqHNi
eiVVbEGW7Qgbtz3B983Ya6o+tsyBCh4IvkPav0u2UD0/eoOdHD88i14jgOF79oZTVvQKvGjr5hF3
Sq/tfLrrL7YBPWLVi4TsuX9qptd4JrmNUamCzhD+w3NdFavJMMibx/9C8DN4XMyxMwbgByWC8+B+
GIyHo4ShosK9kmJ6H8DFrNwC/Jf7+z0Wv0T4mqPZc5qXK/XScSVvG2fGZbRAfdofE33HrcbzO6Vw
Xdl65ZaAQrghBrhf5wzYhnRPIL7426JNhj6pyP5OgKo1jV5GVL4iB7QScASxbHB4rdJhDkG0DzSk
npaKDnLR4cM/ovhFlyuhIo0AE1kRyU8BS98ucAbNkDH+JID1VH9RTgxy/vutwwkEiApWuWlWMiI+
Xax9ihNaNtu/n2O9+RFdv5B11qEjVBFP6X99WYkax6G+0S8NL2pEX2KUE8xAqea5wy+2AOsL6vVm
LESNmFLdrQT6dTZOtHh5ifwcHlOLMnn4/UcCsXK3XqvsIJPPveMbaj6FqI82ZPRJqb99C+cVy1Ax
4MaYWN4hB5NIBxbtb83eCYsBH6Q0JK5zqzd0z+B8v3u98b2FR2MEXnO16r8qSu/w/8Lwyp6zMOq2
46q9p8DNTclq+Z9mgBCBsKC2QFbFgI77XCT2s1x4FGMjv67UO+ktLtZ/OXJU9CXS/IqERNoXkOW9
TEgpdWGkiLGDHnPR7A14NrDOWz/NmelPHlo6XyQrLtnSTH8UAyi8YBL+U4lTCW1Re/jzssk7LSPw
XUoQ2oXJA4eBsEt5DS/aTpUykNkFbQop1cPGW112TfusivpZlnHzNIU8Pc0NUJiAg/narN7PHAJA
HLUa7Pe2sWKsiNEPLWmSyWsFepZbFAF03XVCFPRh5xG2PRiK8AilD3G91o1tBUauF+FsiDSGcjGX
qUuhH0dh1507yI7mAmQlV7ujQKDVbp2oCOUXh2yTq+t4zWqZOEr0F9vkx7kxSN9zAFNMUa1NFa8h
cszRGvkUNkNLdh5aC81ZQrj2jK+igaAf2Lf2lObeWkPHgIbG/BIxZF6SJzPnhjUDlv0jZn/R3j+6
mmWmhBPB7iMuv+nKTBUJIp23s9BRZvVx3M88hHqEm4DlLiR/B5UF0Jc1SbFcEYd4CUPXU/IzwWe3
Fpb8P+h4SeAO2gH7KRiF/PMOgh5sk0JmpCfIPzNCBVOXqSvquIxSzhZqXcw2DLCbGrHcJNvoRtSQ
DWvxX6tgCu0qoBmVTld5dSqQ94w9z59MD1zlIbdOZwUx4flA63gIvjdZhhgEEYv/44OfD/P0qDfG
xB/T1nEtwgMcfnegLcYoMEtNFTOlc4seBwtEfPc5/0999NyE7dhTc9TpkqX2U3q/Lwz/3QURoir/
qGqdmYZGBDZXzGQx2dOfavxOvOSdFCND21ssGjtNeAzm13AThNi2nEPzBl7cWxCUqg0rVE1os1R6
e0j/baQ6SL2vvIiKoD8e1y8jAwWmRxUUG/VbvhtaZUTCb4egZa1VbGWuxEPWwFVZDv5eHq65y8/E
m9L24O8jxVvhAHv7HvsKb0Id3tmt50W2vFjv0jRTKMh3Jm3YljStK1ATA9q+vw7aftt7MdTvMQbE
KSBGGNOXfSePJwiWT2WynjBkyH3flTrE2JIJ3pxiRQps5LbUjT/S6aIhXzCFeCUIWbDOBdWGc/BV
oHlIpO+gi2zyROwzzgAy7UGbZ5FbFMmQo+7Q1w6m77AkyPZLWOJTa73I/PA3QVC+gZjeiCQu2Yh+
XYDnzWtS3fGxPzD/oHOfVhFhYgl+HNB8GK9swikHu1IIWEDIzH8wl8qojPPTrhcxRdF2bp2ej7er
4TufUl8a021uTw4OOcLgqBsM1sfeY390wxqcmRP3nsMm48Ti+dJrYrVpSD2P0P7LBjJk8g76oVTZ
Km7mpAGLhmcPM+oOPMskVd0z3Tl2Td83pMaNkf1HU7jVqlmqVN4w5Xj4B1LbiOl+lDuX4Q3uj18Q
wiibBQQJIvfDcjYVZUmnWi2GyoW5GJp/PJEsOZUbC5Cgvfk0Y+JwgBgWVtdhtzJpbJfsZilDiT08
G6c0YatBHI50HEwnkNtMFcAmwTbd27D3M71iPKn5zYLxl1ipGs784QNlmuZNcKwzFtCvO9YJdUdM
qt0EUdV1Mgnp5RuMBo5IZjyr41ADlTcca4uh0Y/NAJ+THgYiTREnndZ3JsS0g22H2fdZM4+M/yOB
y6qOQs+jKwDi+wQaZO8yFRexIsQHf/4+CJjRUHQmfo4w5Z6Z9pY9gLl4SJwGpwgc1IShRSZY0eXq
29/ig9dC15PKAbGsNKOssyJhFTxYPvCc0gXi67t7hrZViBWlC8ck+7+HOTnoUnBwjwohbt56xiz3
Wg4jPjT4b6Y/W0tCKf7vNFhVswLnKK7UF6kvbJ47jo8es2yQqEq4036uAp/tqwH/5CtF0a+Br9YF
M1cDRgprjSavenKVBze4e+poDjW9KUYVnKO8xlb8rYqjxZGcsiLXkqaIPD6AS54ItkFV+6qD3mZE
orrtpfVVtFMQLzQAp8fr/qks8Gz+Mzao2fV95CQ2QnpDwSA4uQF6+38rQ136A6krsZclHeEC+Yi7
8sWkIK5iztZDGUQlLSevWSbZnMHR/13W2YQxFjl6zMkjX2UPWvpTqPzWm5gmJF4SjHRkiY0ix/CI
jfopX2OD0l+p/VxBNbhV4kD67VR2SZgfFEBwJLcVE6YQOiqiHu41nwO0DD/D7EMRgj2BdpbG0KVU
oTMhsPhya1u+Pt/c7hQtDIja0eRLtlN7UN05RXU85Xd5/OIbVPcsIpeYFYXE6PSRLWUrCo33QgKM
N0paGkC9PQ5wJjaDZ0M4rxqP549Z3X2Ei6nCdg36zRent1YrzHP9T5/81NaoTmuzBSJNZ5I/yBNF
BcXYtMGg1dNXtGYbat0oWTkBbvAsXZiVDyH69RXian2s8UXB74pKHQjbq5K29YrXydkamnaPi1Ep
3S7bcHu4FXYnJ7RBPOAcotDqf1ro20mAoW6c68M2dDza6iDfGLSZO9lfVkX8d70k7QOHh3dDcPZb
vGD2Ho006uNTg1W576yB7BqBQHGG4eqWHnVNAwnSCZZ2WFTJoeIv0mh4+kIWp4dJ9gvw4ybJRwlb
3bbUp8KipCLBTagXSnG1gwoUV5NYUmO201WfYaJok0YNbdmFKKJ8Ar76aobQTYYVs/N3atzPKhEz
9fyW7Ahc4iCxyjzgXqFTerT+MJgpbEbyw++sGsCJW1+BpGndUvQbZh2i0SkrkqKM3bCqx1SJswOP
FjnCJYKbrwNp60HCzL91PauvOo79/FGxyT9tISPOqET1K0fw4AUn8Whemi5cKLx2jQdeTlmqYXZH
YhrUA59uwxDHYo86r06PXVdpCU6++83i7tyhnh8Bohv0DkHWWBqVMXjCQdRBcXX5+DbUir1Y9xFQ
ay4Oov9iChAjmKIXO/glVc+t2tzdOTnZtcPdhqrcQsjhIjvHBN37EU1JVrF+zX+VgM+G8/93swLO
0bUaJA/bViNMV2rFZxDM8d7Gasr4QdL3dtONZy9KsgbItVmIpQ9O1dxmML9wfsIfSt5d4yvX5U8y
W3Ju2W7QkWgFBNLpcmwaksateK3QkrZ/KJ23nyZWVFM26A5MZXuehTW3fID3udkTMwkAnHWhr8sh
cwUMdIvy0emErvZjVvVK09K0OnIfdc7oB7SIfcKsOSEROBdKqUg+6/BTZEw3Z30Wf7Cssek2R0cE
2xYYmL68b12PXBk2QVMJST0Kpr7QLZiL5fhMqE7Xpe0j6NLg8i4/ydnwk+2lj542WUMN691yrZi+
6dLvwxzC8Z2yx3Wfq7Sktw/cYluHA1L9OJSNjNQJdm6SOLYBH0CcoU+KPCLubasIQ7t3XlY/jRsN
zaysJn76rouI9TVH8tmtDdfFYRfXJDHqKM/NINg/DV+YPjd2Wfux1EtPt8QurZFFFqr305ySdh8s
Dc2UwvNuXT+MlVmPKi52KfwlFOxaUgwq2svPl2ienjF8Y9qu8eXFSo1CbkBRbfkDwjgRaCas6+s2
FKsA4HihQnU/gPXuxJ5229kJVALGPpbKovw5tb5eE7YRDqffVJaHGrdThJ2FSNA0i6ZfhR6M/a6N
Ed4yNQQylw8jRSoDrPlVwGaJLnssqAYS42pelkImVgH3U6/IvOBOnZ7rn5h/3Ulyy2/wA6gQ86kk
eTFtIMhyH1SLJXafrXWEzQVxkQSHsodkHBkRLHNWhJf+/I+63gPpezh9hBG1fXs5K+zaAU9P68E8
2OCiHdnPz60Q/g5RXuRa+wgTJTeXXtw58aYnkUNeORojgeCa5l1KHM1bobcjjPsSqgCKbd7jQS3a
VfswHiFJv0noB1YhMGcs86VHvKkyYomrtKmb85OjghRNfZLVEdMfJp1ZpLXltPmfRA9O9WyNJrM4
BfUiY0BNedDT4ATzRdg6IbD9PhcF7Rcoolug0mQa9fucDI9FUmMscr30E3iC1mPj4zSmMjP34p+O
bRyHsv9jaIObUaVDlJ+mZ/OqtJQV7wHoKsoOWmKYveQsQzQKgxgEE0cxVgjKW/X5soOfE+Lii4zf
ECvdRdRrKff7xcdhnfkrkTddNE+8bV+KoOd82r3VUk89mTeg4Z16kAEPvGCniwhWxC5aPo1OFqkT
PDrRtLUJGRQJ2HpcVrKb4HU3cO5bisyGkt8iB7nzKmaHdU3Fvxr5kl3d7m2dWngeMvI5oBtnurYL
0TBT1bQdo6CLWrSsfUxpKialpgVwIb8UAmlweM394SeHYkyPl4YfIxS5wDla9crjLujdRzjQlHcv
TTsUjYxWCy4hmD9IHxKD33DjKJUwVP5R8AvpgMHpY9T6sVsIy4ug22+gAfg9zy4BO1u2K6kzL4Qi
aNyYo8tJLsG2dqpZrmYy2tCAm/3gyuWqJzD811WLGKc6Ai8hkIK0McnRBMORYrxTQkExZOc/4mK7
vbDtm4F5z5shCNBGskeeM602wO07vPwcuJseq4sYF4hj0pqCQ2f84XG7Wk1S5imK4RLDdNhtzKhu
x8o0mpHMvZTY3kyIK/Cmc+mZopz/6nmCrXgqPRRNO535NxQp/J9MY5suHGtGx5zHhwhgNjwpTj6h
FH117CL34w4Re7Mr3TKOqOcmbMjFzeZKzRXOgFPRHaDHAA94btIciw01gkfGoyufBf8Fovld0o3U
ow7dymrCasiXQePivm5E0ezx3PAvKP71CWbi/BuwJHXkaU1hqeLUaLxgbgNjvcxLtOROJv1iCEmp
KazJznwFTCxcA/1inlydNATrXbAEi85grUdhuMAcSvPgfpJxPlq6bP3W+zW+fRPIH5E1JGq2dGoT
TK/O31M+H18fxjT20xeAh8SNP5DRNEYgRWMoQhGn0piO5ND0RdKaJ+qK5R0XJiS4mcbNEfdLZ+BE
l7ghWjqDDbgYVlmfKehqevONXYGYdL1L0jRRPllW4j1aRPETJ7WspuLFsqoxXe6jgUk2QPuhaUZQ
Heh8TgmgVBrjS917bAabFl458f4oJYmlDJ7qJv+iIcnIc0u3b2auI7kDBp9Mu/JglzS6mCKkV5VP
wMzH6aTU6PN6bGu8VQWefyj361P/xB+d79ROij6pxNnmwKlyr0SF5Dj5IuEDuPOZqES+frMBY0Yg
qql+uX43OFPF+oScKmtkV7VxX9rQuv4EfTjDwkz/RDfkCKSp2Vp03Zeww9ofE1vChXZ2uj7Zenj/
vu3AoUPCxXHbEjmYIba2lXliqsxLC6OrgqnhnCgie9Ps3bBPyXOdXer31r5hXmNCAX5bIqoad/x+
z3JLqK6KL8BHA5DDqqY6mpESJwUjiCW+0qCfaj/IbV1Y/Bis+7CVTFemiCpExstcpmAKjzeGIHfx
ArGTb4aSl8PUUjTGnkMKDQCfiwggIln8LR3NrRxutf1zFyz6nos2h2wN7sFH2bC7CqiJv6Bqvp/O
VjGJYNfoI3qRKfaOs/YM8+nN4f77VNJnas9dhwPDdtGCvgWN6oOyIJaDJfHwVSTHoV32O/IMMGyS
x6DzuEYq2VMI4sYn00ZyCrUykxQuN6bDn2fou7cFHLDoMmsezR76jpAnVjeoXp/6pd8d1ClVspIM
l02SSTLMZ61gslc/RlSriEslWYry4kLsKcFqmeswzc10L4GZnbWb+V3ZVBwjvzW3r4/4fXqfGn96
A32Gy3O8667XG9J9arXGqBveV2MrMK9t/UONG5XVtQfQaueSp5G6O3vwDKD+tS85+XCr1eZA6SzI
cjCBaSD0PwFNo8ssTFqQpGdHuFwc+0czg+GnaWN5FRCcm1URKU6NgvTS9i860M89yJ8YPkjYVrr7
9JvWT1AIuiyqF5vTlrORxTzKbFVw2m4SZ296XOWA414T7/rUFL+it7IDykrTuw010nbMvj/sV0sH
Kw77Exw7w7en4maj004xzjsQabii/qNVsEe2L5g07DiM+Vmd0b0HGGP8AdpNBo2ZyiUs4D83ZitZ
TFpaagLluUE94JV+cLDpJ+D4c/FYkrXaEUq74QCeHdobe8uOuj2F8KdBf6nN+k6l+ol6V3C+F02e
5rvS/XntrpOs8mig7cn/VkQXRTlox1UqDfjTHoi/JGFk2HxE/fquiQ8yqs1WPImliKlLHy8JMJU2
F/G96hiV7+yrQovgL9PWCf9HnYZxWcRI8a6uoR8RvHjaOxbrlVrZ7ig7GsUtE1mfmxzaeq9L6uuF
ELEE1MZQUw+dj5GKzmNxsH1gsDwo9IU4IdAVh0AxTZG+QrRtq8jDZVhqYvXvj3TsWcQUeEKm4DQk
QFow4kThJZmOUj59Pwdc6uQKQ5DApC0WCydcH5m+fGPIIcAwmcXprpej9tTH3Ou9Sq80KTp8nYu6
XFUrYc4Z2V8GKU1xg+sG3JQtz56VKMtg3g7OfSXheZPOjp4VP7R9Kkens2npNMQwt6qCGBy81CSH
dOJtpOU6W4mFFJnl+SyPTAXuiOh9Pe5yWVqmZ1pQZqzrz55pKQJCKOHk0ZEFwQU2yNd1JW3JfDnL
TLbRqCN7t9lHL93a/6pkWwZewxR4h5xVPPLUhr55vdtD9vjKl6nsvCdjj5CsiH6mrPqrpj52rr+1
nwVJ+k5gyPIfQG+S2aNr6/uXz0SXFm3vKHENXP4VdLEZa/BVyUKjSUPX7OryldKqOqXI+BC7A1rf
iGbb1oVU+hdzOS9BZ7YOg03Jrne8RR93OFMBSMrV+6ah0A0KPMVrz1i5/SiG76Io+dhRS3pJO9x6
F2KJ0z6tbKNda2O01JAtfmKEPi4kh6qJ1XCK9BtJ/Rzcg9wehNvDIYdatHQRD2w5hpaaxtrViVae
Ah5/lPJ8dcNWm4qzhQCnAJScDB3cVRNvRZKUEczEMsCouIyefAR4uXX6cNPS50uVDfUi+rZtYZsZ
SOcZcT9I8idplNmeH1msOXadoa2cohB1RvYEJFkigqejcfSiDMMRSOY4cLc7WCEK4A7sOis08J/v
Ua/KjcrU4xDlDs8spxHDRWN2fxSX+fsL7A0sKqQIpEiY6P19r2nfeYZIP4XjIA1Xm0y5dTFgqgBE
tDK/J2G5vyR2aI7E+LIlquWLMYKapAZuB8iJHjx7jmJKKp7eiDHQFcX+DIq7kUI1zvDByFXoY1Vb
27cdaHW0h53Tn/BjluNK1cmMBAdGEja7j9fbqFV5p7I35M1ppeFpLaVAGyHBNCn2GnekhE+OGfCu
wd88Llc6L24xU9N3ArR0pUshETmB9c4SCXAEcJAiM3Qshcp9rRIMHJV/OrbFRyOiXV+PZJSfaONC
m1uvYFJWAq8xMGDgNRhiLWDwSMHfjy9CcDrq1fmOt6DkqtPH4AUgtNJdYQDmvEJkdC+RAQYxOQSS
tk7VeBjSyXXgtfef8y+vCcC/CcbDfG8ZxHsBqWeGTkSrjiN5X+L72ne/5S4s1Bdwryom1subpP3q
XO5CN7PJIt20SXA7SrrIn9guLgY9pdRFpXVGZHU+N8JT3k65ne0Bp3bZlKXO6G7b4Z8BCQNj4trr
RDfYhGTPlDqVNtlZdCQhx2OfwoZjoo3hdnK17HAU5dB00qlO1EvKNXQWJGuaIiu2CR4FId+5D9Kp
xq4+ZV3lOM4M0XKuThGrZgz//8Ju5W54CWDAEB5kmkb1uR27s5vVPgWWklXhVDZeZgXUnQgQBJMW
HFtN984FrBoY4iThi+g8xmaLbcCZ6GGWXIBXiVGeIIpt8z7j7d8rRnDoUm8RprTeLdNH0boM5utk
o0ahSM4Kko6XUhfRb5B6D/OGmVzfqy6FwdNXRhm1r15qacw7/L5WwqhucDqEm/PbPwSwkaCKSeux
bxSqbvPuLrhro1Xq2znbWYD6Uj+Z470Sv2dcFYeiBMBeWaZ2jwpnoQCrmUfDCiDRstd7rVDIFSad
ESQt9sMsJXdZEkUs/TMe77WwOe7wYm3zqGzGtuhYIFUEqXQHq3EFEinbaE9nXQtgWs1qg9Xdqclp
js2y5ZDkyOwj+7Im51vnBU9iJ0LGyxyAhrkbD2S+FQGD5U3lKWZhgecn9wYFUGU3E//t7G4UCqGf
pNkOhU9nP0DmgVtAhWHhHqkkf0w/ZT/TB9K5fz7Lo72+RiK0ps6tsAUl4L0vTUyNW5lxSO13ruEd
6YHK8q177voQAMayyCetDvEzWeN1tInHymyModCkhat+m3f0ttZAXSw93vt1AApD53BGiSY+Mbhe
wh3zA+gXBlK1hp83Dipuqg0uv8CE+IHkVYkfBig5vOsOvhSy9i+wvRsBlb5X3OhsAqYwEP3GXOrM
5+d0mTzHMVDPqMZIr/tMfny/wC9UBVVjUYXYfnKQ1ml+0g7DInhdWtOaqukzdVA8hud51pjk3EJL
IVPdLKB5j1r1V6EMF2TNw/SQwsSG5V4JvBEe27kfjKqmPBPN1qc8dfkznfGYQIv8ZuCjhLHvcJbn
K6aocDgfgVOOi7gxxqQbzwpYFf+xdWB9l09C9IDvovD29ZXRY4H+o0IDuCx2yh/krL0txExEfyh9
QVpHVH0UPo+2OzBpmlTdKZlPWCi211FHaNu/cKAZRv4r09NQXI7d0DF2PcOc3KU7LxXJR7E6tSBm
dx37FsSiLL+OMKiWdUeP6vBl3BcFWccp2XoTMiyTfy2CPLJS4rqvksU7x+JaJVGyJqCzDc2PwNW+
8+WJS0qvLBZU7xcYiynclY7EfyDD2BBoltsx7ISH39nD1xBeyq9ywq9NM+6y6euUQhjAWndivA1u
eokwDdmhrTjf8inYnzTtBXj4KIWcw5YQCpIcTQZbuUysEs/S4QAgZf6su/ajV9hvHMLejinOssCR
OWAPb4Z1dVIApudvjtNiVsjNTF5QMUDo4uAbbSfnJothIYyjCoJdq78kqpdeTZS1OjHqfLYgpY9D
5En1ZLHi+cJy+8rLnk9K6Xrcy6OZW61yezjxS4Q5gjmDVCSza+qkNv8coEEHCtmisJr3hOEOu10q
7AuhPSwnVsWBxAnWO3uzjxq9bJOQdWtlPhaCYS9DzbeM29csk+w9G3QLU6OOPeiCESAxoNplC6Sp
DJtNG8KC6RkxkmZq3qVPBMK7p5OFtJHQR3Zp7x6sFTgtnFTCzdAFUrycFHiXU4j3i6bGLShBzf0r
OrYXXzaVBS1mvCYou9vVowR0mWpdEDT9hZlS6m81TSE5i5jGvqsXLaFfgbewiJS/7hYyT3ovooN8
drz0kszV+2vHUEmp6BLenzLJfZjG/LqLZvXCFCexv/9S/AgEYfvOH7Mn4Z4JA6bf8j/xTV4eWOHu
+RvG3EPf7Y4k2EuSVzwKtAf4/r7PMYyTJex9KAxJ8pVNqM5aUwjJ4pq0gbxoRprBwHMqXLNEgtja
UNmoTfMIdJ1ppIAP4edyL8HNB9pmIOU8WR4VjSy1WZ0QBX9WOFyviniYPVCWgfA/d0SJCQSUQBkC
8p/qtnj8hjdJkFmBybXut1mhgL3HjH9Sb4ZJbjW293MFhualH5BnF96snGIqzcgqIWLYwwl+jW71
bU71Aezl8UUytgspFJ+bInpUkoQYIzcS+idcw9uJclElzlvz3P+L0iysYSdv4Ej17ogpzPdrdArj
zFLSbKQl9r2QWPYYSGUHQZXPn6raiaPQzUvNvd7XdFbedWP4tKTXTNYXjGgrsbsI0Fnl21o2u1ec
K84xsHIRvU8IS057vmAfo4gNxrnt4Lj1ppl9XeLJABJ3MmRMEenoUcsGD5Vn99elDBIB37LDwYc6
wD+LX+FSIB/UFQO+F8mAr+BnHeVlg9DLHP7xh/D1ySIKGOoW4mDSi/RxWA3H2mgokhuskcvzEWLi
aiTEa2lv0sZTcSzoka4DY2PeM1T66ODhyKoBBv1WHfMH33ZaikBtBRTkGBqDDeXevkP9DfviXxfS
3AV6Jqyt0gwpySc7MRkOSngNzn/OPqgrODuYTaKBog9wvInqx5l+sGDEgcjxauylpPrQvKHpvjvi
0RU8Asy+3kIZJw0OBflf8doewgFnsuBTdaPJIckCga38Wk7kQAtz+Vgg9IKIKTE0tZxMzyfIALZi
DvN5Zhmmxpu7nD6bfMYFTRdCYUEod+4tzUuG/XlleuFiUQNL9z6gnr9TiUlU0SvsN3sqtg/1a95j
SSHkGLYmh8/vwFpix/ndzIdsFCyvan3jkZjmb5CQ6I9E5dcTGuHo/0XvvSHOnzGmbUEU4+3TswsJ
ZtDqBsXfvZdOzzgkSUc/MHVVif4EUwHSSlW2t1ctHnr7O/Sn3DdxJPJ0BaUoT+EbRtCNxSy44648
7pgzF4mM09HGxd/FYKvnkfak6w3gY7BtGne7biPYkazzj/xCWXJ/CwW2wS+vjfcCe7LuPvYxsDy4
4NTOPhGCsh9A0yuHsCN1sbeJLjJuCu0xTZ+5PXt6wFACjHAMW2QENfq0j4ZCRQ/99M/K1I0UAuo8
yqJ9qtBUT8zYXLLi9YKa1TwxM4tqtDszVuguSRa3FS6/E97rjOv69J3ySTEDtulr5yljibwjun+Y
5XtTvl+DgTMCR4g7gm4LHYYYgj42O3jsTU2IaIJg2dd/7VmNH0Gugm1Q8ZAHt28pdC/+CnnQmPMs
NMt4vp+E5H4DEvxBs4q90x2uGQAkuyagjsH7Fy0BfoeEStLtfgdUpAgzhxNCB5W0VODYyK6tbgzP
Fd0UUhBfzQbHPbojARSy9/wn2iKo407Oh+zpmiQDFVWvBys4FEUrVXSV1qIS8jqdlzbqXmLj/hJQ
YRoFeq+ynT8gqD/SiHNQyG3oFx0cw7eOOAIeMVKF0sly/dFUw0FY4A6LK1XuLRq+Ol8qI7KRXvJR
etOVI5S0BtxGQl2Au90O/OGx5nLBtp1X9zanoIAEw5ICKw1mchv4o5HsWhCXtB0UR7ZILLHEt/pb
WQfyfUn9EY3NVdkSC052MlN1vS7YiwyU88cawgborCauxFA8tVCsXp7scssL2LP3uZ7pGixQsZ5k
xyh2PfxYkjG1vnSdvCmecZ+vtJ4P01HyNmXdfqRdJgp6QbyHjXWo5Rx45MkkZ7CxpK23ckSDabll
HUAH357wyv4uYbFeC0JPzZUC93Ei69YTkbDErQ6lONnQx7lF5hj9d1yF/CdlFju2JQCp8HFlFTlW
hE1aH4Jzhx9BnuBpqdFmUjEg6gieI1JForaCxsfzAnNpddo6ac8pZr/m3etigxTyROzPHMJOY2ar
pW/B1179JHCZAdPRcK3jhGAWhPErSQk2UuYEigoedY5Nurq/OgdNmjNroJmjXyKEmG9UdWE899Ev
iY0Phtlwoe6E85upL0mF62BKaCcviuwOfooBINmiuBLAr/Tch+5eSOgVI0tMYREWGpEsHN2txVCU
fdQ3qD3Hz65j9NPZ6UbIUq0g4Kk2MYNm+LV1t6C+/Eb9MtZSCn41FP1HCA4HKNiG4DPEbYL2Cwra
mjRTBuG6VDLOlcTIC2q2sEZw+YiBfncsJyKg/w41+wfTeSwBr8fSw/p5yKQOfVJmIN/hgSUecpnE
o+qEyB2aBccnfECVPGN9OBQUSrwN2oHo6sUTHoBZwfjfMQjGVitjDIDl+2BkZoya9TS7DAGJ5VDi
9Qu1TeaNZgRw9U6uM4TaQregX0tuZ9F7PZ9yqORnqBNNk497rZCfixQcpRA75z/7dKv2swtQ4Eqj
caKh5eCNJTNMglij0i1vChQY/T6WItxQ0GkxdRA9nblQGV3hHzHWQkCVyhEf6KdqP6C7CfTB1F1x
TkEZ3JNuu8pGBo9G/I6b0gIudUMJJ9pcTGcDmeVIML8jlW9Yl1wBNHlfE6n5seul8hwj60CAZNY4
ZKmUjLL7c4EdBkils6rpVJSrVxoOSJnvB7mjZaZZk1crCt/SYD77W9yru9hezDNrWpSVJEgkUCZg
xHv17LYNQ4b7EVMdkao0n3ZjEkiNKqQCotmjssi66nk5Sv4dc72TbE4fCTHFz0TtbZK0mvMPbWQu
M8o16h8om8rIVBDnS3fKTrZKpfYYJAVEt9AoZlZxyYYacmD0mpANCA+blbpdoduYKiSUEZiy7gir
vxaOHUn4X8X+zT5f+sEXaXvPwWP9+godEc70+5HVH0RKBo7wp+4vRKqyk1OMECSodGkz2UcEj6S7
xzQ3FDPdg/rsecf0HoMktt79M8B9/dwNn0l1s/m61VTTHtH3zRK7lkorggJmp/BmfggGCsdREby4
kA1OrJe9UrKsbvxLWwbtom1mTcFvpBtqtIDqTzcJzP3z21YeQ8LHJE0crc5RUehuy4Gx+RMTTIWG
9UltjyO8nRmvhqdY6OPmmEW+JH34KmePY3SR1+oXrweG3t5WyqaWYRYQnNJvli2zzt8ZOh2frfMN
HTkuj5CSWkTKIrgIrjr4uL7nA2nSAZPF3hKbKs4hvS4CgPCgq9YVPT/kj/3WEvXEdigbnT4k7/g2
xLSP5lny3gHO+gokX7hx3AI16kGaCH1jCIx8A2ulTQJElhnpVWr/izwoYNcbURJ09aPNZ0kyeu5b
zP2TrzOkn1ASfHjalr55wYlAshGF3q8r9d4qjb+k/eK3+Z4Uo+MxjeDp87WhkcLNfpXNYBFBpMdm
JSbftyCTj7q86BYxt9VGtOup5JG2XLt0Hsn4Q/5nveBsSdH/AKfFxaJYDwhde7hoLDS/Xz4uesDS
HsIP7Af++NrUrfK7ZJLhNO7kyLQsQnJ9iXfaZw8c0G6iPhoV/O6NW6BHpnTHUPBhJY4wCqtakmwa
1+Evpb6vMiw5qKXiFv3L4vmhtXHxkFocvgi5VNGb/MMYvHYTasWhtc4/PyRNbM1RfjVdHK+SUpzu
2vxDbfC6VPs2bT4EBH3VVLuMFyexoSAxbOD98GQ4wj3vSb8IygtUXPWBGaWrN6E2eeG4PzOszK6o
dtSRgoG3FCI9Sc+tLvrIFX5IGr2gOMMvZmV1HmDSD4SN9bq48C9/wXMBy34UafUUcIwJriStM1uV
fx3iDb0zTv1hKIw/Y6bSO89Tb9OK/BoDn8Dn5eUmjTlisuhmNz+7IsJrP0/+n1SLDOvTh2J0xgpf
y3wKTVij0Op2ffkpDLK+aEfsVGtRD7ctKyEp3kiS5nXLAAJg9EfJ3AVtuIzQ5G4OSBQ07ODJiUMa
NMIcykGtzdf61dpSc5CjDdqWtpWyPlSyl8cTm66sR5ZGoOxtdvfURrhelrxXZSY8sMUBs/qBT0rM
mXmGcLpsvujZrtGBrrNsiq9MtzwyLBqC4DwKyTQjPI2mbwN8Fgm3e4UWmJSXsKp6rlGXqYmk/9rN
/+wa+bWs6FGLWOz/XgZZn6sRV4EpZh0ESXkRnCWPEiDofnBh2rUL9V6GppvQ2kvNoAkMJXDN9EUQ
ipGBy1z/0mYlf9WysZ7H7NDdEOyK68ZUeztANSPBjHvR7DDT0Gbf9WALNEUMPMi4Atd6qnM1pxYO
iY2UQbZfhhCDc6kO1wjZKVY3EpQiY7KGF6Zw6rWOQK/Y1wFW8hN8xQ0UGhLDOXA3wls13r8KcCm/
AXpO6ZXG0fMFewCJKHQ0oaktopQZHqPtr+lCh5dMHt4mK90aKY+gYjAT/lBbvXnHNtmc+7ksEyzG
jMYidbgNfC07VDISSW0zn+1jVqSST34w2iuYpQena8QbGcIA51y+U3XD+5ABkP6l4drQJNB3xvnc
PBGem6OjQ23Jr7CKcol+Vv+p8rstTXVqcLDdVFk/j6FW0iw9wmgkizdesemGOFlChzzmaHtW+I9y
y671VAhlcuhYCs5Mw17NlJVAnWhUjqxHWR433MvmRr4HBarjLc0Og1sEPdD4s7DYJnvEgdqj2+LQ
UGRjSo9bkc1ErCkBctoVGATBIogVSInua8NJV+dgw1BqvynPvpS5EtksRy3g1A5hgjCzfJicelQd
o3Xsbi7XZue5pDdc243M+x5xjdhWfYw2bRo5B+s1EFS7NBtkl2J8+uwQPAsi67XzEL6RdFor47cM
vFm09vC0p3R6iIhBh+nMqaeQMcmhAYHKKm2+q/Po405Vosnu0KXsmdAccteQ9mBHixIOgFODrFbq
lw971EdY9bSlHE6mbisrQox4dN5KnXQzAw4ul0EYv0jkhBstVk081MX8qJ845vr2nIG8KM83vEZS
y/uHxTZ7Ccr5FKY8Dz9xKM4MWzMFYGqKbvPwkxpxhz16qxeTRIfqxuJvPPh1YD/yzeaccnYxmBLX
u0D9vPnmFeyIT5LUeYeixggZ6adXhgCl8uS23iTalI6Sfd6N4+JjGymyvw6Fc6QYAadQo+oxAj31
TS9sdD/eWXrJt2UXM9XERbONLSdQ4Z9ZDEmKp11/VKFzVuZ/LKRjS4o9MsHpoV/K9qBvNjkIids6
jKMzroNigJ/Vlf8TIdOJeYaK+r6vSt4ZrR3c+xUa5Rb+muyq/KaZDwNThLSbrC9Q/2ET/P7Br/+e
D7xYYmeaNyBoIZjMLBJLwhrDh6yLiZRLytFO6eorLQomnJFtyF5bwHn9/zHtHbQ/1AlFJk1pwNF5
siUQXq0EFUp3tsEunJEXVyAOEn3DHw3nLRvAEQMBmmcWTWoYU4W5Ug0Dh4EN3d0e6xMaCJvnxv48
dAzddQJSzLDhoSYX6PLnq4i++H91iyIX9hdcnXOnImgSB+mYa6AmVac9qGhNVGh/vgrNP4E55H3w
mlsoWByZQCOZemxN0jRQTkP++jcv4NPzTnX971ot36wSQxoiGw5kaKMpHHDycGTnxvUWoHFGa2Qi
0oD1+0h9AoOGKAFqWN8BZuY1rf+b1scs2wqqZ9ExhU8ChXCO1SqqRRAOElshVy4NwhS01A5+cVCQ
8b90N8uw6Z7JCtdqQSmW2d6T0pON7vzS6y03JChXZ525oU0hVrNROOa9sF9Ltdx0iUK8vRNdXH1M
8qVXoaXm0e8+9gdOETkAbZZNUlltFpdjNVE+JGgWq1h7Z/PcjhUhaw4D2u/OK3sVk5/cneTYNyMR
HKjX5jROxCjndSWLZYZBU/+xgStV5GQdVaVii/C9yt+nGRLglH6W1ZyQP/rdopxmOupYm9pr6YLl
VASfX6Ve3hzYqETI6ZgTonSK2SJzZoI1kcBVAyqeYuYN3snsgiV6aHNQEYaLYsLXTEAgsd2C6REF
/QMvAB99kKcdJ8dJlLe9PA52rLYQNasMW7gHDvoUzroZ0RTRzXsfAxj465aFXWHVNIvXIZX3AwJv
V5MESOMvpR07d01wMvFpbQGJXbkJnSu2clHjigvJpxT/1yPcNwjcoysA0bOOcxtWjjXmYIKwXKki
B5MI8FrzVc5B8MVesxzegRnAYEjlddTSTlfdXEUUtwWETB46GmJt3vSjCVt7VHUjnAH3W1bb6oeZ
Q0ZFfGu073eMgvVYVyybzewQr/p8MhLnNCJFFTMhxU+VMbIFNwVWm+yEp2dz7MjxNz4ra8kwd4aj
hOxLXw8MvS36kFyjtxrvwuvMJBAcm6xqaxkCkwSkUtdWXt8Kh8n9FcUXe7t0NywOBfRMUxnCw6mL
WaYW+eNBl4g4Y+9FCfHJGqyNbdEcQ7GhBDcx4tkXEuEMlsGxZwhBMG3S5bkN2D9a1+fy9VFraPil
9Dsu2KDCOhCz1V2tPYU3BzCuSOhaglJqMyx9s+jZTWhbpB2NiQybmZ0lt90iWh1+hF9GNOjz66Cq
zIKRebfwke0S9vlMRJSAz4bOn6s62i8V74VrFqp6iOCHP5tdPTI70/mxxGkMIJoA95/eKeMnlv86
lzMBM60bpssklmzkX6dPiIyETyLngGjns3yU7phRIOpi4T3xPBP2MhWkoltGPGBPF3T8WbIUqgM4
6xZccePHIDEGNCnyLF2nopO/DBN22adcPrnREFFfJ2c+qeIQI1yxFHc7pCjdRabneHr+0vgznClo
opkNUjmF68r/MfEroWU510JuPnsEcRpXwg95Ij6F8O0Fh6u7YdGBCvYnrrHtGpOgefhalFZirmo6
VkcPUYvG/ixgo1Ntx0+JOAZXX4aEoiX+MFypqIyJh9Lj9P6CFL4C4oMA51yqeV0sZ78jHvHr7REW
3es/GglcJfvJwD9iPpWUpVpS6tpkzOjLTu7jLKZ/bc8rX/BFEsnNOzZmPKikmalXvQhDRpwat4KO
ArXtjnF1vhnWbui3FaXKxLbfGU7fw6PE/uP4YNqQ6Lpk3K4qkT7QKLWNb8Cv3mwrGPeOPyXjsq30
/7VQ4V7Q8tDH8B84NyBG4wclfNYlZzDmKONG4u4qkQTwD5VeUzIi3x/hmA5WGFRc2dA+dykGRC+D
FBhNSA/nCgVpgm0oOzRj9/IXszprJ5x/qn2tpA9ixBzXYIZJe8mKZHtom69vC9mY8Gknb8//KVUM
ysUMycXGFch1gYLmtkRG94wWiCJQPA9Vz/T+VQksZb0CZ2rS9tmPFoieFjcpT7ofRRgXP3ZeqQeY
/3561lMRPb7inKWE0CR0yfO858GKTtlAjPY9pKTpeLpB8hZ0TevV5zwGUIID2HuWIaeIBlUhQKTR
nbKdBTZezvvwUas9UUlqoAZByh8SkjJK8sLSZHWdLQo/v8LrEIU9pTDVmxOk2hTas/rM5YJNteK6
cz+sG0ONIVUz2uPFsKIh3zlIkpV7MbCE5ExqtnFEHDDb1MGIvdwoTDYpFfkKwcw7kv7kdfztOJTG
dBsAVqZ9anr19U41IYjLuBif2xNaYNWBlATg6ZC88TTrA+RAhZR3GxrcrlXfDWk+XAztjifoa6zm
3YhY5xogr6V2CVp7bvGdGbf9B1RRnrETHHBWsdR6Z2XQeDsBQzaNa2hNYCtn7GEv9EvlBbyTo3EY
M7i3FhsJNFQ5kjzP+/MKZcDrCEYJZI4mTZftZzN+yseIoJUolwxDrO3Gp9NB3nvqjJCbFOEj6QF3
/ZiEB2kTs7JQdDavPNnXIyG2qidK+ntyPaNoD5xISe+RxIZ1YapmAyFlhUdhsomGMemxlQqT48yn
t0/OnZOUBy+MmUcL9DzExFIGxzje6KTaRzubo77zQxZUtsEKaEp2Fep+vM+gqt21tiDxDK839N+9
93+71BJ2tjk00J5BkdkDm5p1eqdHkBKCr+zZ4yrm8MpV9uDR2WNg06OnR6qtl71spmmHN+FF6W88
qm7DdGkKBLWtYWaXvAjIjZYWq7TVgnZA7CKg+apEyweR7vrgj8yqsRSbeiLK8oxUBag9c+379sk8
p+d8ewLlssqDTns1NaUQgMCantDYlO2Q4iPF5R8QszuB05+DrT4nXQk8xXN0RL0Sq1rFOMKIpvdP
mB7vFh0XCbmH4In3OgXsVRlHxfgN16i/HE5atKhR/2cCEn3079eLjcSsJnsChOE/rR+fZ8rbWonz
dgTuQwVwqS+63Z3f4NKRRHjOULoi/emC5toA8lHKfzeJ0PxD8dMz70oOYQh1hAxY18VTQQ31ADgD
QtQA0EVecVs0vpyOlFvdG02GT+DoAAqRxVCMCccGbb18o8ONUC32bXruBnjPc+K6X8l6FjyogrOQ
9bkM4tojrEdL+nR9a0zcVLKAgVY8UmQo1VKLeAF+3LgkDmDl9C5d5kldb0hDP2zP+KVvrx4jkG3r
LwXVDWDFbnmO6sG5hBZGBsyQ9RUTYqCJZ4JP4zL87e/dn/GfsNJSjBTYLJzypQ9AMg/zSVwqdY4/
8MhmbVPmBCaP/Bqb5TiLClvQ1o9U2hteVfeqRKIN5uDWXcG7zPXxQ3guvdd/uugFZ3Rz7DMaTM5H
vT849H3MVBKcAQaWHtOTBzA8w8onBtlNM6vUcSXuBKUePUnhx314nb5upiuaK7qfu2oeQ8eAEuhY
4PnhLAVhp624+BQS4m4lPIWgE1TPjHrxOhhDn/2aDyxCpLb93pwuVm2LQ2GqDf4hjJwddOXQ2n5d
/b6IaxuBg+zONSGwA8i+Qx4h6SfyXDg+B+oRdarqN4iZb2063quOiv/v3oT2wrsJf9lmDzfeYort
xIP5o0rqoq3IVsAaL0BeS+ldraeMUp3ZEJ+6tUT8tb9RnALp8yIadCejNUkPlREQxydNR5rJgfFA
oF4HKoAS3mKv4eIYkVZamzxviQLOueHapBeK982snmAUukMJshhY14VECbWl1DZyxgxcnTBYFNMK
svy6Avg1j9P0juSiSETG/jHDAN4TV91TcN4erSxdNN445kcv7xOIB1a12Xgr6/71scs3kUaBzyR6
yFtiMeU0SIa+bqSECYpqmsyGvOite/IbO5JdiJjCrTTHGOPelhF7ZP71o7rvXEd4Iqwn3LMJKK01
lP8REE+IJNMq+oVvMi1Pl5SJ9WVwUXfKnSQVaV4FnjNzY0ciobFTa0wMiTeEjy70MmIqF79WOf6i
0SaKZW7IHJmiidu10vvr8GA6dZYU9/ca/wkhmahGt8b11VKEl0Ok5aoKz32XfXyUu7E8Rs9WauLk
jyBBlQue/Uo5SjbsmOCcC7UHVjZ9bJ8Nz+iPo7vIL+Nx1phYq+7ppj+KRFafltQeOAbkRizM8TPa
G/Ka5WGJmC3IoQztuWeXkd6gyDrbFA+L68428e6IZQlGIFBiYBiblprTVulRJUrnTAEXDsRSw7ZK
W5vMFmaSs+DZTZcmy4748eTS8bfhvR+OL9EkntFbRQqPsgptGUNy3LPEPjvwAPmT/mEeZ60A/435
U317CH44xrJrsqosuubqX+Tktot1k/ggJceqEfhkENabMb+puqH+8Su5fDGNuA6RRNeuGz77oJ/y
dG5ooMY35hnvQlFVXFdAbDKq6VZAFv/+9uPRtbmx/MJGQIuYTsC+BlEa0j5JSg7R1kNHZfKQNcdP
laSvMWHYrkGzdmz166LO0K2ZNVsNmfr1a108HDYQ9e0rC74b/DS99/6n+9d4W9fsVVidC+Jbr6oD
0zyxVRPOeWAX383oY9748p0izPtkuJah5qHd8FlHhA1Ddrtv1DYRthpivy80jUX3F5q1TYC7jUPh
jRa65Ko2gKzBPut5JU7X2nae/yC8R8ASsmeTPD8p8GlxlTWWd6SOZkHlcN/3nlDReIUMy/pQRxaD
hnmIyYCrAescbKEYDmPcH1rQeEKOl+G22PoMJ2NZVy3wkMQn68e4zpHakZPVqFLKum0oTyr8VKv0
QKTtDIhRETXXTyemA34keWcJjyuXY3RpbnIaSBA9D4l9lnCeicrt5DYUOe3Vkr+JC7vosEZfAFk8
jQ5HTr+8iT/H9bBPaWHAHjntpfll4aE+jcY9XM5njbHHvxRe9OPCR8o40MBCnL8uEEL4/RHqWZ8g
ufpXZA/HsbXhe9dpJ76iTjwAUelr4Jt0BwU4Fq8EzRqzX8OfYEEfHLUmTTWQBNmio8JTdqC1tm+E
Q72yyNWshxMZu68wgnJCmbZ46CBoMCVv4MMQK7+Kwb2Zq9G4ousIkWmy3X8X2IlRvzNponFKX9Am
opMNqEzF63QMLS2RjC6NAg/aZy4X6bjxfzGu+GmLzqPhMrWCiAkAvdaIZhfhcFwjOXVP2PM0nMyT
QLQOrIxXbtXRsuD6DjOpQuDJ7nzPrpxVkiQjIL1AMv5f+jHaLCygghUadFmBvxZgtNybkD6mjNqh
OGcnbOsqFS185yHqIO5ViFrIkhqiVhYSgt3NbGemqCXHt9Arm+SlIeAk7tbE244j4eSqHYiLeK4l
nONVUeKGmN/aeTDzUrYJ5S1tgQeya0sF6j/RzLLCyJ+hcyQxpEC1KLLTy19NB3zdCIwOyESbp/ve
Xk4BM4clOXTa+ZE9Xl2KvIxVszaUhW8rykFOAr+u86P6V616fQ/JM5kCjNVT7KTgUIPJO3+tc3CV
TKIOccLnRNhldigICNU+TqAeDyioONDiJavMScRJ4g/pT3U5jPh5Q0I+XIQQnPbI4pKHetmboIz5
RlGVvoIkpmyjI2r3fe9WEfzs7KpRR5/bpwRYdRxpb6DfZRmFBLCj3oZ85HLen2xh04lBbKGXVg2D
W07wieXXFp7qYQMiaZht1t5quNlUvXaIm5/qo2CB63QodJYAzesZFc7FYX2Xm/Mk+UfgoF5o0enV
zTqesCSuKlYk7yn9KkosVE1Jlxv8h/lwjS1TP6yPtC3N0l2ViN3XA0daxjvzEbUW58ljFV6XMDZs
uIQqFngpB+8B/u8CULAI7K0r3xUO6Yhh/wXeOuCND1lP1OtmGv8dsfH/LCMx1SGYxXwLKfKfrOEx
okekAi/u6O5DC+t0btihAivCSbU+Mb2U9PYYKi6WJimqdCnDAtZK/VL+dmBTnTX9kZSWUCLfOYxj
oKFj5Pela/WTLxBWsGDq2wNZ2dFR3D/Ef9RXiPxiKIWPTDoG3x8lgubHfRVnxq6sFhP5sd8wqyFv
upU6/h0HsX9sVDwxByz8K/5db8+7h6FL+naKpETceOSk03MXQE8nxaULLARVe4jEdQZu03pW6AKV
ZQCqa2a1XHWjACS91NfpgP40tCip0IlK722X17ojZU2wRKM+LJbPl18ujDI=
`pragma protect end_protected
