// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H^#$^Z,03;$I,K?78@61H?:MPS":#4\O1D<>'!9; 3XQC&2;X@;TTX@  
HD&7,%W3W8L2+5(C4"11F]O3?6H>W^9&V@MW*I"!BD ;#G@X7F)):*@  
HW=Z2K[7$A<QPYT00J5Q 3SZ&+#.QSX5)O,>,P_JWDS6G1&+\-Y_,I@  
HS\AK(AATZNU;[6W?5@KPG)).Q\&U&\Y,MV/?Q'*OTV]E#7%CBY9(S@  
H:]N;7'#7_Y'56R&K_\B&-*:.4WF3&T>_/4!B/ZVV9AJ KC[2S3]P(@  
`pragma protect encoding=(enctype="uuencode",bytes=17904       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@.W5T(]H),C^JYGL_@5^];$?DBPYZQ<%85@1XMT?K](4 
@^0*=OWP7^;]UY7L\?/$I-?L&AU?&,+-IO7)0-*J43O, 
@YM#Z5A+"FI"A-"RY[=>KY5TCLRZ3^J?S[WDUW$*\@2\ 
@B67@N:==Q*4:-HLOOJ#7BM -7K[=S.UQMN.0.!I>@2, 
@"/P. -O4P'"J^9>-LJ/+]H@X+V*F+S(=G[(>%C$/"I4 
@I4-:9]T^_OI?A4))N_N ]Q'SZ+.\@"/WOJT7P::/PGP 
@Y5BS(>G[7/PO/QA AD5U@0&V8MH"A*M1%U,P5AR'+.D 
@UO@+=XSHC-?7-#R3R=+__1#.[LKAHK:#6R\U @C-^0L 
@.%;@Y ^?^.\,0$AE@)=G4-307X]XE+#50A_NF!A>0]D 
@"EU5[51IG,H-2<U)%C(WQ;^7H/S:LWU)18"H[9%MK^, 
@:6C-VD B2:,Z:T*C*V;H G X^]H.C>+*![(R1&B:9.4 
@%?W'X!%R[[CNV)+ 7EF=J^0_XQ .WRP.%"'^IHM_&>H 
@*O-JMCGA5HDTF,!!J4,+@/[EJ>!'3V_]K@SP@"AQ]2$ 
@]84%'VV%9A423[!/P%R[[[&__YTWUKVBH8#MP19ZJ#X 
@SHO?!^4S\FUJK**+UT180;UP  !$C0W!&@480\'HZG0 
@$)XR3;&0EDO75I!T3<_A.RY<M,+-+WKI?H194)09:?T 
@/2^//G,GCH-MP@21/U1MMU51U%-B:JLC!#N&X6%N&3X 
@6DF5H7Z/O3$L,F01,Z8T]J T;=#3O:^,9VX.W>.ENK4 
@9,J#AJ/\$D<HGFVJ<2V0D18@9\U_V6T0W;*\ZRZR6KH 
@ 3V;W^*#"MC>H_*_7J&>I,?692%-H@ R^^LZ*$/B3DH 
@JCJJ;BPA#D4-NF@8I02B3.V=0?2S:NG..=.]RBKG+2< 
@Y!U8N A!.LI7F:9*-GB4Q4A-44ZKKHVH1XR'+IYTE?< 
@*2B7KX5W 3I"Y;J=;L6/WGQAA"NB<#<,[<_) C0QQ P 
@DS[N'87[KF#(CPFI;=UW6IF^>P7>V39.4+#]!IS_#FX 
@A;WC#OR97N2JN]70+SV%H,8A@1%@IS5.0 K&C<B*!>$ 
@DM1P)J8LM;S=X6@QGV'3U15Z!$!(#\V^ZV8]"+P/7KP 
@<2YO$"AG^"T*! X,CI?=B<<(\5PKRJ&G:RXI;^+/^6T 
@;[C!C*^/+F%7B)?I"H_92R2_M' 8"5#(D5<=E_4V R$ 
@6=M!^;X%.3(J8<NQ9(0EV7ZX]1.K$G?3)M@9'X TY\  
@G@6^5HS>E+3#A]&\1>N6K_G:0$SFX#JMO0U>=6E)0&$ 
@,Y3Q\FQ2B8QG]GJO0D&R"F<^<&(P!-9[\?!B4DWF9[0 
@K_ML MH>SJ-0G98K$9)?=V\MF,B/A0RR]GB45:(X)FT 
@@TJ;"Q6IH,_J\7.LS0\ZVQ5' L-/'37T6:X4*D]\=XH 
@_TX*Y,.,T__ IR35P%[707 FXRUQ.%7-(SAE4@A/9 \ 
@WKGO'_+F_ORXO_1?9EN]O](23KN;DJB;LU\8A-']3=T 
@+1CH(-Q$BO@=+[+)USUYD,YF5!!7_@[IF5S0 X2(DU8 
@B$#8PB^D>CYY(Z)<XB;;,.PAM=/%)80Y%>*VQ7#SB_L 
@K7NWDOJ,9K:!6WJD)'%SJ5+P?>-4VE31BU9=WGG-O\H 
@:L,<U\E E %E?]2HO3N_SJ5^?/3^0]),:(P[ENVWJB0 
@).'4"AP0<!T-OQ$<;$!% 3$"X5IV^<+NN4G#?G"ET@( 
@, Z97]>*NWK=O$OCV[13%=_TZ*\BN&4WQRBQR]:3(O8 
@4FD(J<(9DDX@QZG");FHBY9O</CEGLA[R+2(CLK#H 4 
@:]NWE HV',! ACJT):_%UIYU/*73\>X(S($-,IQ4JH0 
@C3KN2K1>0-::6D+E6B_3Y\8SVZ89ZH'(84=X"A]0&A8 
@21@<^9DWJ:O&3KLZD=N;L<Y8SO=')=?"RF]7587&0D0 
@7B%C4"5R.T-AA^YR*ZDZ3Q#+X)]_KJ0D?]:B=4[+YU0 
@& YG<F5S,HB$=#@E9!H@=.^W8401_BWW(XLF>17Y& 8 
@7F#>U-5=_T!9X\L'_JRG^?P<$[IEA@,>S9Z68.<ZP2, 
@.;T=D>Y@U]'_1?2'\1\U69^;9/P&ZZOAUD"?JW(('.< 
@Z%(I1]( 4;CWMC!!5,/XIJ*Y\M4D2G0R#MJF?\?(<Z4 
@\3TQ^]B+[*$_R;SF]L)<&X[1R8\"AL/L/+HDT'4KUTT 
@V;>@=S+@ S\+>Q>#+>/=B1DOALY/[Q? <B?BOH(^6CL 
@<?FHRNX0T: ,LXS6ZZ?#2>\P")9VK&F"@5?9_Q_Y-&P 
@MBYR%T77&/>JE/0*4Q*5>L".X9KS8I"G-/X=4:L-Z\, 
@R7"0]7#5D0$H^@*:T0]'N$(TW%/>XY<,*OO&6"2A,/X 
@ OLLQ%!\B65%U V(=&R\049WS,5<CNEL'K'_;9;HJ+@ 
@4J;_<X09M\+L'*PYSSU0@\;E94ZDI:,P1L(]$L@ZI9$ 
@CH!0?DV9O])]*0"4 F#'2AW*) _OEL:)F\:VI5[W5J4 
@.^7<$J3&%(D$?*X^MSTT';U[^FX_G):(;O\6<+O=(S$ 
@S[*@YFTD[8C%/&UV3SK^_"J\5]%$(R6;\/Q?U_MZR>H 
@TGKW8SH"CO7, &+5';#==N>,_H3(/IZ")#$5/-\MB!  
@:AHF>^+!XLG4[7R\67>WO,P!/@W/!LENF!(_#&JO4*X 
@G8H6SBR)UFBSU;(_)!.!I .8<>^'0MD3I&&B>6"/.Y< 
@:SPXL&\4#;":K.9@TB9HBZU^;R[,>,>QG-^[T<4QS?\ 
@9=186 W&^*WRS5$\%W6+M/IV\39H2"WF6%N;8;<RJT\ 
@$"7"U,Q Y(E MC;EX3_I004Z;HJ1GU3/*!M\5)DZDP( 
@?:\ P/QVWQ1E91/R&?O%$+T9'%;P:"4@%6Q^=-98\PD 
@;/!+=(L TWM)*&HO<G8@"*BI*]A,24SDT>77(JB/E9, 
@SV<2PF ..CQV/=7),HZ\.F"W6O["]:]>ORE))F C23H 
@DG* \&2F$M\!BOY3617I)?E 1Y?Y)BY?A$&:BWW65:X 
@UV\^C%J,=.XPGD*V=TLMXD]MMV3YEAVU7Y$K$KV<8>L 
@9O5.B#&Z2UT@OU361@JRFJ9C/A,&V;OC)CH;S <TCE8 
@JM?PLZ[B0MP1.]X=US>M G-\6&3B(4"-&X\.9<E@\_$ 
@+/+@QTQYF-A8""M^G8A+6C]-@7_3 O+&K64<&+36U0T 
@R02,<(?1G+.)C & YT(X7"FJWFNE[S23YS^ESH0JKOX 
@YH <G<LNRQR59ODP"I;F[Y85IZ]H/8;/(;"^I"FY>H\ 
@+098_&3)GC]?\*-C"[!V3:#2^ CY1KR^8L=5P&98_K, 
@!!?FUMHA,% KMLC^U@1?*"ISSI7'][G2.I>>S8$.BS@ 
@RI0-Z(&8B'O;?C(F["3*B@NI!V*!RNI 4$(V41NH4=4 
@SI/<#XGOQ5Y#J9*T4)%WOVD%9)I4>PBG*V0G58AA %P 
@Q<Y^IA1!"2*H#=Z^!*.E_WZL@]&70M8JEIF=M_Y 3 X 
@F_=[0HIA4L9[]F]YZVA@D-+'H(6FT*%#@YC:,HST4.P 
@GR*V6!%#HIL60<]"4^V'&'O?&B$H'!.IH\E2ISQ@+>$ 
@DS*@-K@ N0(/6Y4V[W4!=(KH&J>SKOE+*?E:&)7N^F4 
@B;S60[A'0=*%1@KU*&">'P@<<R/.K6Z3 *36Y.C7H4< 
@CXQ06S6)!5;G&6)&;=$JW7(M*M6J(QPB9F1Y]/QIV"P 
@''>(%$"Y=GQ;'7E6YY@(92^ "'L(KC+NG]RQI)@W%Z  
@<,([B;K72\'9Q3F2D0'!-8 /ZS =B3]ICJ>6Y",(-UX 
@-^C^7#SAMD:'Z_08SPDRF?Z@13F'H=T;G:X7L2HPTIT 
@XIB(/;CR9"]70] M'6NM5AG0.U=(;IE-K9A==^9/Y/< 
@#GI3TRZ\=\(S;+[-\/<7<*WXDG!CW0??7;QI;QUE9\L 
@@5'7[Q&8ERP]R;KJ)*'K^/V_I'AX7YR!=*?#2C1S&E4 
@."XD6+#1:!$@+AALWL4>P/-,U'PX!/V]?3MQ45;U4M@ 
@4$D^@_,SYP):VW?K?,C'WPU>W(:>3\O]^''EUVCL')( 
@OL,;$/6UGA#6H4L OM97&,$9K8:GD,4B48Q-:TTL6F\ 
@6D![5Y.JF=^Q62U+]P=D!N?Z;)2IWA?5<-%.%IK8'[, 
@VLG4/KR6C<*=U96[RJVBC0)0(T??9#V4?ZW)1B;+8'X 
@^*2^=/V \,A0D6_UPZR3$-(8QE^"R7JH+I(B/+.;O ( 
@2KY )$6+#E?'6$' DX=KJJ;M+$>/QP9$">D?1!(LI%\ 
@.27<!W^(H<L,<PA)R BDJ?I,EV^H"8OQN,.EPF@<!_\ 
@C ,2RU?L^.93]E4X?CGEX%5DD4H5@$!;K1+ N5I6"NH 
@[JT.*6UN))2/0(&E58\@XOFU]5.Y<CZ'.WZZ7V3 &-8 
@ER?76E')T7# &\M\>4EC-O6@3P>\&1R>VJV3IE<JFJ0 
@T^GUUMGUZ)A7[@/R[C>Q!T68QRGBG-"D2K W)OT&WJP 
@T7^@1]07WFI+<,>510+6$S%4[_DB800J#D;6<7F3VLX 
@K_L$Z3<C_=)#VXL6]W ?FG"+6UG4<V>M$-1"L]5X0W< 
@^5K@K621*$-A@.7/]".J]$FY]!T-V4H0V7V6+,VL$MP 
@");4*%VJ_H_>:GC5S&4:"A*"%(F9/16UFV*T&"/P[U$ 
@36@>J7"&4I].PI)IFWBYPC42LY/2X'MC#AR=,0*(PHX 
@B",1:VT\4ELNEX%[W)SIWRA;"QU"C8QZ4A4]"\_UP 8 
@?69[3ZX 5JE-*['86#Y6-0>;-O=X?3QF*G/W%TCX@ND 
@QYIO\D8HE_?]&<2YF,B7!$^6*<K0N/5-U5:::NOK#\4 
@,:,A48MZ)W/?]8?..9='TOLKZ(]N^_#T F7"<*>CQ%\ 
@T8UDMI>R4N OCYJ"U!MJV57% J9\+'3 DHOCYG87J#4 
@UOQEQN8U_;OPFKL$5I]X _ 6+K2W2$VOJ97<76W\$[0 
@;=02MU4%GS6W4A!LYINR+F\XR>O,\E;=(KP4?<\<B.L 
@?F)W(]E4GM4#U:^\Z("99?'L(^N['^I;QG17JS*2Y&0 
@]">;4?F^.L)U^2AHV16K@H3WHI./:B8S&NG"U0>_2T4 
@M(;HK&ZFA@A1$C]@AE\HZ#=))A%&F==4Z!&37"<L1]8 
@5BN:)-L"17N$N3I_G^.;%C^S?%JO8*OY<[O2\TVWO>P 
@&C<8@+14R=,'>*PL3V,@,MHXERZ"^IZ4T,(?YXY 2N( 
@4SVDPM.NN5$7+&2_#6-E64'!*'D<V\B/)IS(Z!K&C3X 
@K!R#FHW_C^AY7#^=TJFQ[C%#<&^QN9[(T9R][50XC^H 
@1-Q'?NK-H46N-7BN/(.(ZB:*;;)<\48"_PKZ!-^-DUP 
@#BKR+[_]%>I+;+*;SP71@ 7]_KVRR/+ZT2S=&G-Q>9, 
@CUN6Z@G@31#_IS2B8]R\-\8+/;7KK7LL"%T1YQ_-/1( 
@;S_H5YSHD3?6YQSB+SC[6*4E 47<KOKM;C( $HM<O   
@(Q6G_"P!]Q">-X:]LC= FLL;OK.6RT95G=A@;PJ$O^D 
@D5IIS&\POH4-;>H?.N22*8+@N,#X2A"BK^QDILO<T=X 
@XFCU^0LC"-D8$T4@<.)Y(C!C9_EX_@6@+!Z;(*-+V1P 
@_+;RZ:<$HW$&\W6-@X_%K" 3!.<H$'WC8_ $Q=G;!LH 
@#Q&@^&[B%8\T0'XV";LL4VF?3H_"]#.HT<32,^,J<<, 
@6OHP\1Y?-R!@=H _J]B8$3B5##$,H!.>VF^)5YQ(#L@ 
@$=LOBUYI3=896A6VNO#ZO:.JJM_YW4_ ?"?Y\3+,) H 
@_P2U%%8 N&R,<1&N5WR"6[HJ$"9Y<C*Y[_9OV9?7D.P 
@<*'?=^[Z:8;@ZV,8CSNA=9+AL,,I?HPP#[X*\Q_R4H\ 
@=#%Z?AJCX,VPE@?3:+9"-/WF/]P/GBI>CS#"N-W%J8$ 
@= 5+B56O]J+1U/"8[;!#T(/R=$QEA3LR\.FH"JV:P1\ 
@M)!?_K8?*YCEMZZ%OZQC<#"U[_B*B^/F[4!446WEI1D 
@['^-W]R6SB*=7SN:PO,7^(3#XD)#=K%>COE3TND=EDP 
@(P&M+[(.3\E(ULADC-"4%[_-!V_?P3*Z#?S65FNO;JL 
@*!%K_, _TLW^?F<D$^./04)L5U#6^+_?:*,4FYNL 9, 
@O7.XWJY9<[*S%9Q0]N]KTI<+)0M3ZQ-.:Z^^/DW+J'$ 
@Z:-P.+I+RZ[A*'*^0Y+N-?5MRGRG$U6;1O.%-(0VL!@ 
@I-'];N3-3\0_6'YVWW/,VHPKC/\ ;C+G)WHD4L_0B0$ 
@WZV"I1U:L7>W?27+)4D_*%QH"($Y)U>)#A]\_"XE'!  
@L)-JL"<LMQNWN<IQF ;PL#<)'WH6;(JG78H6%2<PB$P 
@78B]DUG,$9!JTQ&<UB0Y<"T;B&_&2)[B/M$(6Y<OY%4 
@$!3Z[GC<2*E:\>&3'FC0=;>,-D)2.#+%GPYF/@M/7/8 
@G,*+#G-R^Z"_H'&&;7H)&>RWP1#ZWX_R-0T0W;I9BP0 
@H2PM9MN*2/4W,LJT&82<#O5:T; \?EEAB7AQTDO;I@< 
@1>'.HOMB)?KLQT69[&_>R4].1C\E]O53;&[S\"0,T@X 
@/T&.<J=I&@K<PT@("YQ[.]4*@ !=H4&!X].,Q4:M"50 
@D__8FY1.<8A-ITRP<<,4.B4D\0]UE#&ZBE/F29;/(@D 
@$,;T]!VS:1A7OZ1R_L^S/2N*1]_?$F!NP+Q"]?.*N7P 
@R,.>$&;3"XP3+_F9Y[,C >R 3!"8&P\-->=SI'QZNOP 
@\"8.WC8HR[KG]U"MYA37OT?,!%%,9)1UL@IL2^#<-$( 
@OZ7A^;[:3&<Y[>;MK.5C6NB)0U" 6Z\<UZX:@]NE,\T 
@*2(;EHWM:I!PDB\&)XQ2B,!;]/U50H[ 8%:H((XN^&4 
@9_-^J 92 \(VV]Y(2S5[ACX+_1T9^;+U#07R?/2T#JT 
@&@M^)G.T%3*&JB?V;:NDXSHP>#/H"#0(=0LP&R,'@O, 
@J$AW?"6,5'&<!^'F! E+=P%!SE>6.:?M>$D'QRCXX;8 
@N"^R,AFL7]1^K_[#YLZ(>J0YA?'Q=E>-\@4H\C*@#>D 
@#M S+*:WT$%R<L@=+Q[@JLT$W908HL&AV_IEVB7N:38 
@W*.RYPL3VS/#0]]VJO@QH%\D3#LW@;$*!G[F:<#.*[8 
@IL5,E0W_M?GHO\=")/^(: WIKGK@6?<BLKPE5Z<_O9X 
@QDE(<Y>.[:10#%&4(V8:_)Y)(/%K1-,'0AV#H'!%'-0 
@Z,!CG?_BQ/K5QL/[BE4:]AR"O-.L%'/&7ER@E@ZN*R@ 
@@*/Z3"""\MYXE3M\<\11Z2\L9L:W4LTPMN(V9SI^*U  
@JFYR^'RS[[>M_=GV5@#%R2/0SZ&DK<*0P-0;@9#S$\P 
@) (I?)45YD,2TX,$:VC?>Y.;!)=66N J+02&U<QK!#L 
@*!]QZC(>@(6^HL62:F69>4^#1#:U US'FKQ;Q=V,1'0 
@:'_?7;:TH)KS[&-KCU/Q,Y):(BN\Z6SPPTM'*\K57<, 
@$R]2MD';H3!-@:IVDRYK("L3:AY?OY4AR\9_P-3:IO, 
@OJN+PM)&JC,OSE4[+82RH\#=\6X@JQ(R!.A_#T6"QO$ 
@A5U]%G/F;:&_/[W(;7+)TAM)U( \AEV]OSN8GA%7O$, 
@]&P(Q>=&#L$Y[Y5U,%$*<0P]_%R2']H4ER9^0F9YOL@ 
@M^ZN;H?U92K:VD%J#FEAMPS1J8G%YD"7-V+7X8I<#H8 
@L*. SC)#X?LWL1#RZ79%MW52!\QZ$3,]$*!4G]*ZI0T 
@K+H%I#[*O3]+/EF:0U$<1K1A+T1.&6Q2,@RD\=E/C=  
@4VC37NY22N/4LG7S\#(.=+TJ3P2Z5J/,= CI3#Y& $X 
@2//^V9>G:.NT[<\8#AK=>DT6?"]]P%P)]=O2O)4%1+T 
@I_6M=8<;$GL_J^Q,G+)8@9N<,KL4?3E8;S./#+>@]ZD 
@V.D('9C5,U? $_8G.\GB#>B^#C75)E+P2Y2H:W@!YR\ 
@^;N?N-<G+92<J]U4EW ^P7.K&CLBR*>).*=<<&&=6VH 
@IK5II]T[5/^^-.G.:.8SCD]48*GT35M((G4BBNR23@@ 
@.QZU1JHO[]9E'**)$-6!N(RR"9U0A\6?+FE<(4O,-2T 
@PRRZ/>IKR=Z&A6HMV:7A]GL1\ D#B20B.BS[2L0[V"  
@$FSLW1$5%8Z?!E@LT5C9F;Z/+Y:>ZCLK"D;QN<^THB0 
@)6RR5W^B<B@\1K%">XACZ3V/&X[[$):71I71@K YU], 
@'ZH33OD,>Y#&Q3^32E$,UN#N$XA0+7L3O_"D+T.!V$T 
@K1$)D"#=E]?0P1'&F694EIK>V#?Y6")7])Q%LGI9'.0 
@H?S9")5KKOP [U4$12/R]!(RA-/V@:*O,SPLRWYM89< 
@N!?"51TD/QJM;<]@4%1)&Y>DB*E+U8T Q==8?#H@0J8 
@8,I-(JYP\^:S-R4O"@4BAFJ,N2YQW?SI.8IHCXM"#,4 
@7V>']M(F+H5B72?L4 LX/T0]TFSNH2KX5PBY$J7ZCG@ 
@\SO)P@@N\Q<L7WO I'-NV!EE2MMN,R5[0I39?;BK:($ 
@77A1*!7+SJ%\.1M_ [Y7JL1E)E!J<7H'-Q"M#V/G8*8 
@-L<.;AA?@!#.$@%=.!M(@]@LCBZYR+G*V6V)_.?,2.X 
@?N]FD1BW^#:]M!42J>"!S5@$]_MVZ&^I,%0?U*=*&<L 
@X&6?UEECO4&E=JM/ FJ4%JCP>$[7MD+]U7>!=PQ/X>$ 
@T 9XE-ESQ<$O8-RUM!9WI4B#X654:@+WE6B#EK%)3XH 
@:X2^YZ38P."[!^\Z"NJ7D1'_BIG31N:4"L/!R2S<#ST 
@N$EMCFI^B]]I>\E90C_.>B8\3?X;5BBW@C,2B<\\&W  
@'*.=V:PMFKQT75TA35>#(9:<!DBCGZXCL<G%4.)DZI  
@)P^0@1RUAV\ G>U*.<T PA"N)8\[WR\X]$R&,*FJ.O( 
@!]<@S./=I7CV<P4WT)MYL!)X%'8T3&]RS,_D46&%NLP 
@O;/"BE- &^J@F[1/6#7$C/APH%A_A7V$\&]Z8&G0R$8 
@-[<E]J'&UJJW6F0"[CJ;[*V0?LKHFX96$S0>9A](3%, 
@0G9BF!%\*-W@##YF>PYVA!UA$PC&\M63-UD4@I]D@'( 
@# U$[WE*UB;30.'G8YFZFX#SO^,'B=]_\-A5_9XV=JX 
@S6$8MUL@&L.,IXB,!  9BV\(QM-BP1[/CU?RGZ!1#_$ 
@LE7ADP,[2#.:!'T$-\ZTM=XTT2!+)T9G@S#0_]>)$W$ 
@#.:)_(/@"<:&7F7CX%JRIY--.922):(QZ#-\JA%<>'  
@];=L]:TA9W82LP1N-'KV5S)Z>DKX@/$Z5#_>X/^=UEH 
@2*U/R#OOTQ8$/0?TZWS9)G-=,$=>=<%( IV>-&*X9>< 
@)G1>GC#^+51V.KGK1;]@SBJ0EZV8%)_+RZ/1VX80K"D 
@=%2R@6?8IFM$IT,7AP+,$B0:BQC1Z(Y403:LEWD3ZJD 
@I;G.O)%O\>/N9=4]_\GE4BK?W9G"0.HN4_?E"6+4(]0 
@Q>+E1X6;>_6ZI]'2U2G[U7$G>)%ZR?2Z3<;>RPT75?( 
@1$U^7)Z VZS2@798:U:2?O$_N0-B$?\6\J/;10KA.\P 
@]6EEBWF6B*\07K=5E)AW.C^"M[%MKF7R5H:TGI#NY?H 
@=EFLMU4W*3A'GI )YR5F<G*7#5AL0\G+\H_>$0I2.#, 
@6JK\^^57+#/!+=;!^5!;"^2 UFK'J-D<0GQX+])>Z%0 
@E.R):>(!.O[9&E&1L2\D8K;)49-\A94@R]5>?3XN274 
@8EU\G%+5<&16\+SC\?#<]LO4^6MV<SE2(#E-_DD(854 
@VOB&S:#!35>+IW8*65G0JXG[XY('<%QC(;O4JF1G/.D 
@W/4"DI1,/_-FXHUI9EXZ[]3&:%//X-3!TGO#=]D,Z&@ 
@IQU[A;\%CTG\:<6C3B<<9YP%[ KP8&Q%92[V%\_9R,< 
@GI<MN\'Z:MZ^W-X8Y,C8-CY=J=!DOE7W#6CN%5D'Y&( 
@NAOP4XC3U;EU^Q#(JLF8;0@I^=/#E1*FK\IOH7499FT 
@=E#9/AG8,3A1/0.O?KD"\J@<[V'RZJV"__N&HK5P8Y, 
@QT^BM>74PZ_-O\EMM(>MUS5EE;='^*,0JTH;DI90P3D 
@OTX3P4=4C@TDGW4ZLQ> @H^F#'G,1AL$N #ITY=)_)0 
@QSRX#-7V%NTXH2011'-7G"KFM(5Z /TI>1("K6I$<_T 
@&/*4.WJEZK( T0+BM[YL3->,1N!S)V!\N*:[>\((SF< 
@/3U?% D1;K#IBO:,@ZFW(E/R=/\,Q<RYM4'6NZB7#I0 
@#FL\CMM?)[=KP*49,IO?>&]^-KGVICP$[+UP&/=B B, 
@.QO%Y/(NO!6@]-U"H$+4RKD)U_!;/*6N?_\"H"'+]\@ 
@F+X]O8X;-SN*\UD2'MKG:]*./7^;U:QMD_+4[\<RKRH 
@7KA[DP>1IZ.1],=[U7^9T]M_G!/8UM:NF["AS5C^U&, 
@#\Q3[F'[#B5PH^C2^TX.QK&8(G(4.JJ^]"$'XE:2ES  
@"^S9N7>M 4Y\.XATP"7DN=T*S4TH%X&5D+Q_E.AEQQT 
@I7%IK2['^-3-&QPT_6(3Q/?3%1)KN1'\-PA <5QG\CP 
@=XV#:"FES/70Z]W0L)>U9\01SUE#O]C"1(U3V"'<N,$ 
@2 4:_'H]&R*=IK"=A7=N/"-/;S@-MMM7G'H& '$*)AP 
@'#@P1B=R$HFOZF3;_^\.J<2&D)^'7&V4Z8O@]7_<+34 
@!2V;FZK-%:'\(JT X%53SZ&;02!2L)&!VY&=CP6 *MD 
@9T[GH2S.X/FFR2-4W[MZJ0*AF>WNF*/4^!/W" K[HTH 
@7=1M@E9&;<Q8#7=*9+&S.%6(<@%N)!FH@] T):GI 9( 
@H^N*UIU+ HACGB0RCW46&4IW:K\@!LFA5]4OT.QK^>< 
@XUXO:(4- *HHDVRR?)^JM)>#86]4K6L2@H[4)_2+-BH 
@//=A%ZI5]M(^/&?,Z2C2[2Q>&H>TPGT&?WM.&QDT.6@ 
@@H_!&%2-I:72&=:LC=CP-S%$]/HR5U- 9_!6OUT'GE8 
@2)SK7:1UN_1!1O??T9:<!K:( 2O4#FS*X/AN6"F:<R  
@_(:#D7'YK-;"#@E_.?5P(]I58OE3I+1JUCM(@=X,^5( 
@K3ZWXQ_"/?1T]L,3T. /5W'?^AB %,7#7@?@HBS.K%0 
@;I1"1ONH1B8<FBX/\V9$W^$#<\_]V;BOSR)[42=E=C8 
@OJ<:E;(U)QA\LA(EZ'5EMMW*B#SCX1G2"VWLX#8<(#, 
@$#ILBJ[_+S<6FY9.$V 34QV:Y-( $**$C!#+$1W*?Q  
@$ *"*!IMU;QLG*^#PH36CEVA[RT5UW@.WV@Y73>)XSH 
@[+_3%YPPK5;9MR5:7'FHMBU3]L65-:ZV[:H-Y!SYV[  
@G-Y?_>PC[+YK!HEZ7[<#*!-0_>7^<K7KP6]%&'Y,[1H 
@S5Q1DS\#J5HR.W$60TOE%LRY^_L!UB'$WR@_SDR<Z"L 
@!-]P"FEF0P8M&(G*/1O>,)-23PBI6$"U3XXF,VV]B?H 
@O]8XQV([2<4+9T;4AL^)D>QWQ/L?3HG 1Y3W9NF8D4P 
@$D&[,D[EUR)Z#UGZ:L&0;9:EK*%1671FRFD=1MV'G&H 
@D"M!L=LPG:0K !V#E+.F 47I:TDX*(Z5@$"7C[C4E/P 
@]6E?/N&1%@TUN_B)D:HLVP8^&OZ!5<(*>T-VV-5$/\L 
@I/X U4Q#3+LS#_FR84)1D9!!98QAK?'%SU)I7?FT,&4 
@=D?X@%Q;,(U;' 0V)QE[;FB*)>-_R(\CP-ZD"&WTIFD 
@3ZQ1#PNHR:P;P2Y,_"TU_DF3@JU0,>_R#[0(UP5/B-( 
@4)Y>N5R]=_QU#I <MX&_J\1;VPW)U]*[PH&FL.@,N"$ 
@0)U9O@^,J>)_"&:?F/3*?)!\8^<:'F&^/ $"L0(NRX\ 
@TN-E?)+"$0<Q*^M#XF0#)S^,MYN]7_ F"PIZX^*F^;\ 
@AKM"?2?M#  6-Q'^J,<5D&5%NH_MQ;B71K_P1@"HX-P 
@66KUJAU"HNG H*/M JO4%D+Z'0H'0K[D#K+B>J0[?Z< 
@<NV-'=?GKE"GY.QVKX+7D>?HE4I:=IR1H>I[-AI_K<X 
@R!\9Z6W.?9.\N-)3"YJJ0(HY=2W<L1X\M(X4 MMH!OL 
@.M$/'WI+Q,%OF1C&\40JTF$TS2*D\O(!# +#VCGDXDD 
@Z3:2+>8V$NOZF/45(+C0+5W4.?5BU/OZ$"-D7D3CW<( 
@=DX&E$;.8BE_7,94%1ZL(>QV,[Z4I'ETT>S')1R[2GX 
@S1NOY;>KIJ43J?9X/AA38-4WAW&4],+C&*9AI89R $X 
@#%/T[RH>T;MFA7UJ%#$7_!*<A-5I2S;B;CF0"@[,Q>P 
@#]XA; RG6/G17[Y&&Q XL?T92]8XQY2-AW]0C(R4IPD 
@H0D_353CG_.L-C&_7S%7.9K-_47ML0M]K-H-&, 7EC$ 
@\@RG)$E8*0OFT@0[=6_3;-WBWJ+,!LU,:V-+6?3Q&0X 
@'\>MKSZ4KD\2)AO0>I K56+CQ33K1SW@3#_T:=1NF+L 
@DC8)V;# /]_?UY6O*[&$X'NUH2+&H4YG@:TU4-./+W$ 
@*3-0T.C6A7]["S'A%/3N#ZS9KF1Z4=7DCN\=7'[$0UX 
@<W**W;.3^J]9F/DC#$ %I()I;"RJ_FV\4/FL;+4C 5  
@QL'G@2QX :;Y/15/_W:L3\)*"X>UJ5_0&$X=B["_]&  
@$@&"5MBVU]1R3(5SU3Z@B%N<.4[E!>UVBTT>FO1,<'D 
@W2\ I2W49*]-H,1J"A'%BF![DI9P40F!96$9$D:3.N\ 
@.6U.NWF$*5Q3(_+RMR%JGUKV.TO":T0<0L6/5IAG^+$ 
@[=NLR,=WL%'\0,VO8*A$VU G1EN]U>IM<FG[_1NIDT@ 
@7"]<<SX9',BBYFRGOY^NLSY9>D^,;-:_C;)ET+/G@-< 
@L7I$*E;!8/:&=U1^UP#$S!M[YW4='F.G*HJ2#H\B]*T 
@9[ Y03*$12;W_?7KHG<5X+NW]CR9^C[0Z-MWV_2*9W0 
@OJ*5;'NLEZ##!/6U$FU@_\:&'8 ;TWX9542YP9Z&U,T 
@)G$,CWC9<&STT\N'CFVP;3,#D,.@T6JZ[B.:Q1TJIFL 
@81LHO7(A<#_:$A3,O&T.L"H0$LT\K!2;37.'Q!'BF94 
@E7(ACAL@$2&U3_-G=5&.D)Y-&",^F>J[EDS"L[#8 5H 
@2OZ(@:NA6#MD.W^KI0*GL+G7W836Z>S/V<+9D)+4/3\ 
@GB^+20NQQ6(*.5,6A^4G6G=1/IV!QYP#0(K-3?X =U\ 
@92,<\)51@L(B/%'M#1;!TFM=#9-9W"-!+9279K7G,DD 
@$6K7V7!PF#^B)G02!>MV8(B(EBV;%!,S" Y<D\"XPB( 
@E*Y[[JX)]87H<J%,(+OI55"7!(K"T,Z]8::.0F50L:H 
@C% )D7884M%S+[GB$;X412Z^BS0V+[4JFU'M;PO\HZ$ 
@:G#">&N,8VQ3(>&B<^O!^\DM-V[HP.F)[('/'^LLOR( 
@QFLO&C)<@O.CU)<=<.GW)DT!_-!/A\5OS7)NC3,V6M0 
@F-^$!+ZKY(V<NV&(*.8<$4 5/D7!SV5Q:U5:)#AHI#X 
@@MEQ]H[!U!4LW=_/@NR24YYHI;7:J#W:UZZ1RN]Q(,@ 
@3G56N$V)FSPD/Y*I*=RCI_OST7&1&S9KC0RKVP40B5  
@,I!## Q>$>NQYK$'._CB5>O586Z<Y+P\5E#&MC;HVFT 
@L.\CPVIZ[B>\68XPE"RXIH/ARNII$HB474OS^@ST;1L 
@<1C$#TDZN8VFQ%'8N]$73MM@F-1@M,P>3(AIL/AL9@\ 
@Y0?EXC]\[H!?^;V%]C>)\0+="U9+;PM%#U=51P8CWX$ 
@ZH7L-X,2YU(F+967!T@0LKSU"?>;G]]'35PM6+LB '@ 
@*9(I5",([\VDO^<N$Y6S2(Q^QL,3&UQB69/+?]A,==8 
@F\*NQ&3QJ+O_YMH]8V?7?48;N\8G*@X4!Z>[A:;@[Q( 
@0 @<M3@@?_FJKH0;FC&PH-GHKICS]ZP<F)$ALT"/F?\ 
@]1[B6;<"$*RA#)3H"MU3@AX/84]L*5$R7W47'C583;T 
@C6X])%%*"HD02ZT_.-D*31@9)B2'0JYXF8ZVRA+Z<;, 
@%*TDJJE5GB==*)V$8RP 1)XCR2\R(F8>]?Y2@*=2NX\ 
@+2N-/$M/79MP/SH%^Y15XGVK9+TMO6+>A^\A07!+%U8 
@0$[+\<_>3G$$?"%A6-DF([V36=U0<>M\T;M_9VL;+'  
@J#UF<YE'HP>Q^S*7EF3'HJNNV9AVU;-,[.9"5J&@7:X 
@;X$JF=('.;?W D_&N+B1^LRK]4;,-ID9/P>B5D=6+ 0 
@;SN5%8X&HA.4*J<[[X(\13?G?[+\B'Q%:\-9R?OND5, 
@^^("Z82SSA")Y.%!@D2CY:#HG_*$WE_N<I;61O_"CU0 
@\B/8LVSUB0EO*N K=;;8LCGRU<3R8@><<7,5\](M>*, 
@"3 A/9E L8[V2#XLNGBFX7%L[H<]FOAZ\#*+83^M$\@ 
@:*,?KCG"LO#)1X$/Y(!^G$PL9JY!<];<M:3UK>QV!B( 
@U&"3:)XFWL9_5^CD4V5\L=+Y1YK(- YB,7AS>QY2H1, 
@@&#Y43_$3+W5WS? 3.S>8/*0K 4X.\G R&GXSDF9 ?( 
@ T(/,5Z'2;ZVK"MO:L.L20\2.0F"6RUVCSUG@/B>SA, 
@@ 6!,/1IIJ;)NH"W& _4D2>,2N+_HSM*8#/;/KT SWD 
@/*32QN'04Z8GQ*3D!C(9LN_F6_G$Y6=W=,SD*L:O"P0 
@X$5Q#5,6]7M;.3P8%CUM*FK!%9JSHWW=Z8F2_+R'PX4 
@,\^EC=U,K,BB&-4U=E# DQ&:>,(>:J=;VI?<XOCY5#  
@)$,AH,%FG7_B8$>?9DB^.2^7.2^7>,6\UA)/7TE8=MP 
@0FE@D/9(4%-';#F4V>?5'WH:[D-NG(.[2SZ2]<\:2JP 
@3K[LA#?PRHC%DT28"L_7\ N$IPW)(.XQ;#'X0;G)9C8 
@$Q?#P@ D/^8SR W?JSA,DT]_?-L/'M ^7N@F;D9EE#4 
@"AA,AI1,]<L:*F)U DPXAL_Y3"Z=J1I3BVU_7?A^?RD 
@69D'HWMY%^$M%4?.=(GY2?N(H ZP6D]J_;3>A82BSE, 
@K7M>L17#P&CPQ^=QF$<P=81%0G#=G3TDGLOFF\3 G(, 
@L,MCU@$B!,B[E)BJ=I/5UG"J'6Q@<-\M(4+3""LIX#D 
@;@"H!I1K'@-V)F2\>BMOR5>ET+4]XL&8;]TM?EH5,7X 
@[!_,UTAJNP#)E,RV;PI@E\M!)%X3T]"WQ6-[Z\:+RT@ 
@B\B5S!X\PKP[+GM:5$E'><QPBR_-VC=9[.$\\>CJ#   
@HDCRL:25N5>;3<5/6CF=/'Y7"X0=,1*0T1NCTW;GFSL 
@56@%ZD4O(@=NXM#7FL(SZ1F758EY8 \('!1KLD!9R)P 
@QDB#G?LV7%TE%+X7W25=L*@>!,P"P?]X)S%(8H3@7>  
@KO:B"\*6<O>G6:#U M \YI(-E5C6_]+EH7KH<5\&6(  
@&BN4=T9PE\UN+5M#JK(2B?\QZC/V!?P )/)G(#/\I0@ 
@Y '!WA5--)\RU.Z.P?Q"&=[@QJXR/?D*)'(<UU5RQO\ 
@M_54#D.] !T9L:-PU9FYAI.E1PA6929^7GR8N(#>/ 4 
@?()W=P F[ED\;U]2]E\Z#ZPZ!UOA_^K #BG^R)U>[%4 
@=@(TD?[60V;R0*%S-@^E8@%1@,5ZA#E#W ZQIC4XB'X 
@524U./? _&KS*4Z"0UVSH*CM-T(A&7K,AD]VN%7EK(( 
@)]^+_PV.B<0QH$K- ><(^Y,6.)8>'8HB ?3?20ECE^\ 
@V0! P87VU"ZPUEX.JD7&(* /-IFB&BU9M4G-WN)&&"X 
@/E"[TGPCY/#DT5%V-5ZN'+<.P30*-Z\OV)RJZ!&2X/X 
@MSPU=[*V -X:V;1A>A79;ODE&)]#,2'7<9G;.\X(>?, 
@C,(] )Q!&LTK,\,*.K.1(%R_SZ]J?3AW+GJ%?+@P:PD 
@T0G-3!_^$Z,9I?D0AD2I-@YC(-^YWI"KFQXWH[_!ZOT 
@,";FCWYHPMF]*V.A$6G%RWK5TE634[W[?D:0OK5-?Z4 
@W/3V,&= '@IZM=@3L?4>:']?TZ9J(5.RD"5'@\O<W"  
@?=%C1WQ".S9B)$)P^H]1,A*QZHZ>1%$RS0KH*^D32:< 
@*4<^>UQ"9H3YH&06(1OVXFE-U%%D8MFE^MBPDI*]:A$ 
@8WEX&/ECS,=*=7-$@5YCX\<J_W*%-*-$KD*132CK!5@ 
@N^INTNNVQ\*BW0KYL?'7V:PMZC*2J5UM:%<QY&N+%F( 
@#V>"[O%!@&^YX4U\L"XZ7REX2D]Z=^>>B%N)E467*(X 
@(CR+LL1;8HP1WM Q&6*WSK4T-H6,8;$G8E.C%XY_Y]L 
@B6>L&4:">1BK?+L]BCR(K%M[ZT?ETMWF].]-[/::=IL 
@]@FL7A\$&DW"F  IT(BLE,,!!D?L?Q QKO8YB%[$35X 
@@3L:F<3'63Z_CO3,>0B-XS%*Z[8APV/B( )1-LG!J^( 
@*8K>E6XV>%,Y5;6:W&:WO#]A!)([T:#->^_CP*%?8;\ 
@I77'+2*I>/<RN^,M1L#"Y*H:LE@Q*L+<V'#QG_-?B9H 
@"2^-#[BZ/8;<9NND1Y73WNM/,V7[P1!P J\3;^Q7%J  
@Q>NF ZRQY95V;-A8,0_XJ"0<)22LUN57%WGNC"GU5'< 
@GLCMVE<789W[;R=U*L" X^&S\H;H[+\CN,N#Q=ZDR8$ 
@%6@E9KWJX+MWBWIP?6LC92N%,2M&I!+0D#&1:[Z?T*T 
@RBB= -*%^P"F/ $^G2Z%XPKLS<3Y62R%MCOJBP"&S80 
@B!Q%9MGU_!S!*+C04R;.D,?$F/< @,<.C%UZ]4K6?N4 
@2FI_;7:A$NBL5@3%8P2\P>H1L08<P**-;)O  C)B OP 
@#85WC6<TM*M[VH2_MK2L;(3SBTX=)_Y=WG-4XB<:J[8 
@N=I]L\%<Y^N'7J4%'?3JV?5D>: "&DWBOGAS+_:);6< 
@Q.> O[NJT6.:RC'D87X2?0K/=^,096J&X2"4I7J&3T4 
@C]85P!DA8%KV"D-Z.2=CEB.80%,FD>T!>5;<3].9@0( 
@<H\C$E).#\H@D(0L;<ZJ!-[(//E?_Z1*5B!<RWXQ$7  
@B ?;S%')PWOR$4>::F['7B0P2@CB+J*9$(-'3Y\-MY( 
@:\$LVAQ.<0.L7J%RZW9#[/B*>(F#]MV.7T"(=&,4!JD 
@&C:J*18L$87=4\0'0>6: K3&HP=?+ANE1=,Y@>89GD@ 
@E8G2IEAW_Y04)<_^((M:Y(U<I+=%[2<-P6<[&ZTI]ET 
@;_#=F.G&P'-3SM]A^9!7XZ(8,T\^$>O%,ZKM+',?_F( 
@M;+0#9C,U*&[]91-!J4HR]BM<R_IVQJ#\I ,?898Q<$ 
@W3ED?>R<^%<-=M#@W5!Q.(.A:KFD+K\5"B8_0$B10!< 
@M]Z=@N5=F79ZUE&6XPV/D;/-6172,WP JX8";SG3*J\ 
@W7\E+PR)5ZNYG[ND1$W"G/VK;TK=A*:UK[).^UJP_LH 
@W-_&6UZ]48(+).;I&RP1?(NN/8)$X!Y ZS9GNT[KMAH 
@(I]#])6&@W&_L6(Y>]B@:?H.H]L"N@,_] 5Y1FLM!#P 
@#CMS2 8Z!;V]/W=@^2273GYT6 4[1S,)$CO0GVR6&UT 
@%[9V6K0&15"_N@U&(#TT H>?IIT'EV!; %N]6F&#!E( 
@Y92&_Y-?#3L7N&R! F7-D4'<3P$84VZD:>=PK'F^ C< 
@^01![9^DRTAO5Y)NHS;,8@7Q4S%Q!3MG0!KE:RHJR=( 
@XP!+\XM-)NIV(LC7WM1BY:BPF5ZXGA!9S!5YR)!'I]( 
@VD9?TA0P8M@\+O,E[ESUD%A]X4#30LW-0=G0M]V&W9L 
@3@T=-DZ=0IB,1&C4Y9SCI0)-$E7^#LH<[0JU$C01[(X 
@3PPWP4#*A$<^M/E[CN9QKL8.,FT"T::?W]ZT/_2,8\L 
@8(0B)3\K<%U0[$O=,UTW -(FR=G+3UPAT_)WE%RT0J  
@ 9$J<N!/-?Q3U([%F R17(GS>1@U8W7<[=T.HI.H>8H 
@6%524>3W_%@JL*UQ/63;Z!_GKR^!.#8MS[>ZEX:M)T8 
@T..LJL[4&EY1EV@T-5\">4 OEC5);,LDCH*8Q!3TF,P 
@&UU:5UI](F0 C")J)51IZ(PEQ-4EBUAU,Z4<2MZE<FL 
@6XFO7T2\%8CR8OSZCJ>-$39^Q^[-/@C=JWI/'[I+OL< 
@?H;J;WDW@OK*LV?JD[YGRG:885+,PZW-3*R"L-)>YY8 
@==_E\Y293;BSD-YDYP:UQ2W<>A<Y%@3ANT:;G5V"/L\ 
@!!FQV[C29 U!KML,]\,[/*DV*Q6Y75Y_Y8/(8;2UD[, 
@C =*R*$D9BX<AE]E'KI8.VVBD!AX;F0K0A "G4&4UEL 
@X%KP8K"M7,056%Q^=Z,A"-FRXRW8.+>_'?A0/[T40H  
@E66VO^\92;.#]+W:G>L>8P>_<\]@&%'9:[&[.Y $8]8 
@L/U'=4'P*%J@ (=8+*93Z[137P_(4PM9A^.J(M?FJH< 
@PA5L66T!H*UAHI[\JZG01R>D'\SO7!/MA6V+I7]<5M< 
@5D%*PNAV05]3X5ZUT9U"?D1<:4!$9]UB+2[X['@4F4@ 
@)0S<U*D\EZ/#L[(U128C3PN?004^^26"5)EZQT8[:%, 
@LY+U?<Q4#[F!H&N3RS@"=(]*!'^9L$^\01.ODZ)U2ND 
@VFMLZ.YZD'S%V@!4AS@=BJH4;[+^RQ@'D;5DP\L3-U@ 
@^$>?5$R-\IV#\U23Q[\%DM7JR>M<".V\>YL%A3&S8JH 
@B@-/+6YK9U'6]XQO#MD>M08X/C@-IL/(.51Q/< @?4< 
@V1Z7.Q!PS &A_4)B,RTW^9EK>!T/JI<R<C_<PX0:*TD 
@&607#ZU5#[YSA3PPN]O6W*"S_R=[2IE3_/19D&TK4>4 
@^U[/:78J&E<P!GZ85K'S'(E!0'#^<3,4#EK&;+06PKH 
@"LE1:7Y]=2D4^Y5S*YG!P_HTLXC477T>GO8UC>ZWLAH 
@G;TPX-P/SA.*P25 M$62S(\RK J=4$)P!\C_\@09[,@ 
@+VJ-<=9:LW5),=L\M2B@3$W<+=W.P\8%K)?I1^GD2<, 
@%.&0ER?D\/W':IH7/D\,R3'7@GGKP5LVV?1QY1/.7J\ 
@8<5EDU+I.UKX)V^%^^=!4#$M;[FOI$.OS*-2V^HG'*, 
@M7+#GJY3G#2OE<>.%W!6S+7QXE:Q:SHYBN2QK4B6^C( 
@#2X^(/]B+);[T<&P_:D8LCE- A8JNB7R%8&AW^@";64 
@X,,&8CLVDE XQ(_&W$HAMR THRO@=YBQ 8[@"W[Z5AX 
@0BRR?M_1L$U:!D[0)C0;[4K";^Y68OI=AA:C(ASOZ6H 
@9P6:OL]_FI<FS2M8GR[12WWGG$D0SP<1M;SWQ_;I,S@ 
@8 GD_C2@EI3J)%'S6H>:$1^NLH,SXC:59=,YC.(;^W@ 
@(H'_ZWJQHYV;_JUSBZ!CP06+!<E,%WH#RZRJ.#V$!4\ 
@V\_EE.@XV8)*_C'>3>.UZ%R(D9U\"FDMH<3BYM$00F( 
@#'[C0ZP(D.#7+BJ)89NAX9?9<?:J9FCO-N&[RA[0\BT 
@A,3HU</^;23\BT;#DATD7S$?M6M/.TII^T%:L:O-KT0 
@0E(O:*7+\3I&JR1>0U^_K0X%'^D3+5L$_.R.G ]_>4T 
@HCR\13T^1L$/U!J_RP=]1N8-".;LR\T;8(-^B6=:3A0 
@1FW@ IAY^AA)CT^-E4 +IG?S,"P\L]=ZOCE;,!%EYEH 
@_.B?^&D\PWRR/:P09H083@]%'8K;ZK^0P=!E* T^.$$ 
@O"A:W9_?>ST8ONCYJ/DR22US7SDW@%LU^\R"_C'P!;D 
@?G&*_>Z;= @A_Q43+M/.B",9[$SC3";!OX$%,/CKN;@ 
@V;B\PUXH)UU==0DJLW+KK+;(W"4<LCEM,YR>_O72]Q8 
@]SR]6O:_"T,=,42BUT+^C^.P.:5_MS$MF'R+BK+<\WL 
@?'; "&UV-4+G_8B>2PE+XEX1%*C+2.SZJ!5Y 4+OKN  
@//B]?[A7B; N1Z[OX(509DDP(E#)NQ /LDIXV''88*8 
@!#<R\<5-;UU[391CJA#!I'P0*_3N[UKFR"@.E]/"C3H 
@EQ+C-1>8DBP9EU ,E?LI2(@J_OEQS$;32871K?X,&GP 
@C;\S'._.+F'\;YGF'I="L+VQL4#P[#4[\>C]C,J@VH, 
@)[$4F'SI_<];F?CY]E^=?"V*1_<5H9H\7G%O7A"O;<  
@2SLWGLUNG4.%7<BID5-#WII")^,P:#.=;.(3AN('KTD 
@J<. FMYW2QLW'=)@B 6%Y^M@'WFNP$>W?!/Q#7,4AG8 
@GT?79'@7!@;AJ/T.?F@R"<7$+7:R/#:*2+LH.'I$B.X 
@*:0I$6/! +'=P:;6&N=N*O*62(<].="!-5*(UK$R]'T 
@# R8HMXK<W+%CD'0UN:D]DF[C!; J)V5R%<IF'9B  4 
@N'1#J'N44RLJ_<)/JCO^$6VU&L<ENJZ#0G+$@T5N=?P 
@#$,!E!J>HV3N]0;C,(R/2T> YA>Q=!(TJPL1)#3<[BT 
@"5&>H)4.WN$/<P >IL95K@/H1E),3R(\Y;8'EY!@/I4 
@E.(L!3+?H65UX7LC0(/A6ZE#RIO1?)W;2Z"FO^7V5*P 
@F8(\=X426)>;7E2CHXR$! S:N@_+W8J;X<4DU^99!#L 
@JPAR$O<C7>3(Q!8S_[^ G_6]LW$?T@/$G%^=I^+51!  
@>M]X-/&E)K,\-QQ4ZC8M+K,U$<O:/"J0 B#']^Y_G   
@[I*1Q^_-Y8EB2CM%S&;\%>_&\+S&19-UN9:)UL!SU\< 
@%OHO3,1W 70V4Q;-ZN?WQCY;7^DE6GQS:#VI5UCZ'.  
@9"CAM@)(<((IEB/+^325"P/S0I.'^SEUQ60['C )G>0 
@)EOT3Y[D*0AXQ!<)4IKYY(->)$_2-E:/!T$"NJA#4XT 
@DK0/FC=4Q&=)4\OL U8Y!7]_W:\3,[Q"AA')3O/H28, 
@YKC/O\RJR^WMM2JT>)9F5-2Z2F+)3BO4$EJ>])44'7@ 
@L8*EX&35Z;_S"9S9WRJWD803B<T5]A&NUK"*@=RIHZX 
@:1?<&VQ7Z$E>R]='0%6+JNBQN,ICMY?"LZ)!%C"AS;< 
@4 H P&S8U%8F9!R$ZXHU8TZECEK/5AHC;!<.Z2W)69H 
@FKX#(?6)?IK#AV!+#!@ ]FHNJ)A@##Y+!#2+_[@HV$4 
@(ZAO1PIUT[\TK&+AJ-=N9\ F4ND@7DT55:YOML>3IPH 
@78J3.*&TJ&] *]+/HU^;S-^5B_&LC&L:M2E9'MFWJYP 
@I(.,'&]-CY4!Y)[@6VKU&LZT?Y/RJ&7*:J%Q[;:K@X\ 
@YM *"IY-#?4PM,@87NUB["EV]?+X^[7Q*)_6?ME$5A\ 
@U#$:"R:!^V#!TFN'()5;DTXB5HAI;!U\P4RIM8>HL-\ 
@JPMXR@%([NO*>UQ<-<83F-4#Z2XLH7GMJC!D.!:?=R8 
@!" ;+506>*UE$N$0\6T$*3C2B3,:G'Y%5%XO4Z.;_*P 
@Y;8WM?8QW&0,Y>POPTV'6Q;QVE>W5*42ODJYRK9B;7H 
@G C7ZS)LM^LZ1W5%EF88#$_!D':;F[D6"4V\+U51;YP 
@Q@4LN :_,TY&VVL0K55OPWW)A\RHVW\+D-J]T#J^<D  
@ADL XE8N,>4W"!1')5@8P)XD)$="$[B7W:**IY3(]?0 
@EV5<C;T;R5NX96726S:ZSG@U/)9\'_3CN- 28$.$P/T 
@7?SZTIGF/:_97&_#@G.EQ8AE]@F2FX'P-09KO>WI_2, 
@(9=-D7X-10O32YEA1.;4,YMU?=RHQ5E@/"]W=OMU'9@ 
@#6+@@/;4) 3^GD5HKI.=OT\C\*1.]A^1+-;;F#.<A=8 
@T/?IVTQ@.(IAX6Q3\M**271X78E9K5<JV=% U^H72YL 
@A6'G@CTB?BT"LZCQB*S-/A+*GSBP;3%KO$Q?P=O:A_D 
@NM3_KNLDS>\I!0RQLZYX[1X*V.:TF]W0EGT"5 N0;N, 
@NK*/Q:/V*;SK@")\?5@>+%H"Y/+RLK%=0-2='1A%6;0 
@_3Y#L'1MM&Q0HF5[ 5N#S)!TFSVM9G,^N/3G!L!_CH4 
@.CF'M$2 U/(9V1M.MY9J>W)\6<('$O6S%)^)MKY47FX 
@8H$7FUSESK:YS83+G0!]TC(<9X@N0)B;H8*YB$_UE.\ 
@<7!^^**8)X\H')P)JZ7_&IMD@\>+90B(\/&/F"(79X0 
@%VP]5ZQK+LR@Y9+>-I[[H(<[0'NE7]'INBOK',.Q6/@ 
@W;/YZ-^=&RQFTW'%DIV]>Z8A==GO@[[1&4^$XV(F.W8 
@7]G>.M(^1*F9(-5$5<>=T@%05M:TDD&8.BQ*0@Q,%.P 
@77'TBOKL[I[Z-)D/5_"1S7^3I7C*.K,.(K"FVA:J2[\ 
@K9  .E;F&&8:,BRF4CW'"UL($>X&Q7-#5]F\)4C[Y+L 
@>%^>>@5=Q&NUNG=8E@6Q2C&"UWPS<AEC^)FOW2,NMYD 
@XJY\N;BD,N)SCG=4 9:W"@[:V_7YZIJ7)W2VLO'AHRT 
@M3UIZ,NYDSVZ2W0P/?W :M^_%36]5 IZ:=J,^?U;B=$ 
@&T@[#=B3_DW8K"S-3W%AW[8)X085,U2?YH9MPBA4^#X 
@7R9S^?(D)V ]Q"\7W-#_"5I1[%QM\E=E%6(44PJ$*GP 
@$G/?^OKNS^23;>>4_1 P8[HE .8AU+&8$PN)BB.[\>$ 
@U"6O4CMMO9Y5AT'*MV4TK2&GL:3&?\C(I'.JD.3->T, 
@3]C422L814A,L5EYZGSWWL*S:P"4M@,#IN79U8TK;7$ 
@)Y:J$&-)D'!WYH,(EM-N%78T9;*_[!=D\!HZ87,7X'$ 
@CDLKI<LOE'+UB-WCS'2@Z/3H:AGXHF?TA">F1/.GWA$ 
@\-U)8G8UG\62E_H;1_Q)PY9&TU'W[W&U6M:N7#DW<DT 
@"^3(4DT/ $EX5!%POU<S3)+M]]O*E;7H#"\-6='L/R( 
@%)[)WXTCBAQMP/9UWHIL&A$2P'$&O^8+D8;A5U>:O44 
@/F]$6?:#Z]\ %# Y]\V[$0N.$KD?.@R5/DPKQ<"?JP< 
@W_(\Q!$I KAXW !]!(7B#H92^7TLUQT*[Z#MFTDUB\\ 
@>1[-\/)IB2!KE]!BE#C5[2N;4]&8?!E&Q\-RN8TLTF$ 
@QK;.V-U*<TY/"-R9K>>?S1MA&(>_;M2&-AKZ;#>PE)4 
@2CDJ%%UJ4D>;YQ9Z%L6)@XI2UJ_-(GD0:F<VQ6$^VWP 
@(QK'"\\2"&$]T:,[?BA4-*F*KT[N&'$[M- .+PM!-!@ 
@0382*D2K,M9AYD:Q9Y1N0-CNC0+<*G\_Q0<\XC'.S^< 
@2XB\KO8?5(@3(PWLMA'SE=E:A_NFHP X@\[&3QWJ#X0 
@"G<RV7.6;S^4";%T875TG#A")ICP(H+(7!>J9LZ]HO< 
@G<?+($:"NH'Q#**2ND?3S>1S.AP7KK$/<<]3QR)I;#8 
@1BOUM<[YSADF6)_$H#%XST_O)G3&N%JI5=*>LM(?[>\ 
@U94MV:U%G2']H[ 2Z9B(:R$NCI]+>! >Z+;\?*AQ=M  
@;F*WDUM*"H993A0QX[9-XH17,8BBE\>SQ(<_3ITL?[H 
@3:AM%6Y*O[+,[GS*)ZWU9>!/RL2'&ZR[X'HC:<EVXLD 
@Z(P(S]0[Q*]I\]1OQJ:A'E5EGREH:M5MV42GG<Q@06  
@<#RNW1=<_$#R__^2.< T/F?>X&H%R-DES/\O>@;ES(X 
@:I49XTF.)%$Q8RD[P/E%R6P ,H,%KOFFNL.56"4U<!D 
@=\\N.H(V)B1++C% (S+20B--2SIBB.)O35RLRH$JDD8 
@/$YY41K,2WH=,+SG6;!_SS2X84.ZV;%L +*1#CC]H:( 
@UCM3+ZG5V>T3,PX+T<8O! Q\:4\P_6BP]VW_5F/#+/D 
@5\3F80E$  .UC7(]T1!O3X7.>.#R7#F&F <\@JQ/*TH 
@",#@U-'P:?;3R:>CX2LMD:&V63+:!F+WX672@,Y[H.\ 
@?,T*LF_&>@TW"I][<@F>%F/9H&Z3?6A UM6] #\A.1  
@@J&YK,FMH-69%A'3QU4MR$M_\\56";L*!<(BJ CLJSH 
@.*N79%RB%S?SG.'L?*G)/JD _E]#-J10Y(14>&AS=V8 
@:==&Y$ZTTFW)]07TC-ZN=XYWP?V\K_K$Y!D?.5X_/V@ 
@PJIE?E[C2W5+>.X9F GKQ@'#OPZ'K="F*H8G01T:Y $ 
@1\16\Y>WP^"7.^&,,GS _#(.3BZ?5BB)R)Z0J"O'TJP 
@TE7+LN^-N=[&;\ 1:0@82PXS*9V0Z?FJ7:&3D'1$/V< 
@#:3*A*S8O).9J!3MD.+K?RV;;%\OYC<#A8<IBGF#"SL 
@9<;<V-&BK/=.8S,"X%.TC]O+)-Z6:J0>#[F,B(9U.5P 
@9OZ:#C-LYG,"/H'D!%B/H**"LVY \14;?X*?&LB76O4 
0 JAY 48$:(3X.]3X53[QOP  
`pragma protect end_protected
