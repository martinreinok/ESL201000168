��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�d wr����)S��G`�vY/����tt�V6�!Ƚ�^����IA�D66u��'�-H��~Rhf��5f����,�y��1i*~�
�M��.ի���l�gUV��o����4�3( �ۇ�L�2w��h�vo�/.-S�RO��k�F#��M&��&�d�!�1	�^�AD������z �PD�A��� 	�
nr+�i�7K?W��G�	NIo�(�AiP�_�Fe�]���FRӌ �WY�����(M�����;�N~�]�K��nw�f��a��h��J��9����>��,Ha���b�kl�FՀ��]�(�^�H�v.��n���w
b-!L�Bk�@�Úf����zr�d��嵞V���bP���jR��� <�/�!�H��7?B�i��ɀ;�V�萝�v��i�Rn��~���L�
���$)�6�yƿӒ�rnE�ƞh=�kT�L�����]C�qٸ!���߭��4'1xՕ�XRݔk�	�	_ 2g�D4 o�߬�C�X�',S��.�[�����������%v�U�e�ߗ}ˀ�MO�Lw�?�!joO�M��>|��a�z�����i�&1�l��em.&aQpJ�J�����ј$�Ef�&Ji�?����7��|���E_Ȅ�Kdq�X��/��6<
B�3���5@���j���s"�A�G�n�RF�0A�B-���iH�[I3k�l��<\���儳7���/�g�I˖VШ=��.�|��AIA�dx��{�<�v?3����?X�,eaCUb ��\��D�#	�㽿|�b�������;v?f�>l*��|���MW���}�����]�n�x9��M4�V:��4�ߩb�z�8yw(��öhh1�����!]��;E�p;�>$^�~���0�;}����F�~�8�T!���܌켼�ظ���|*�Lao�M�eh�2�]���$^��������C_�K����V�gjX\�xSi��+][F�Qw���Pc�DF)��+D��øUT�&���ً6h����B������_�/��8�M�S���TѪ��]1i��S��!� ��+~��dK;�FI�v:k�а��Nn��))(x౗��!�4_0/PM��$����67����)NS~��
�F��k?���x������mf)�|�a�Y[\�u*��x�哈aWu������e�:���TI�j.f��^&�]I2̶�����o�������D,Lz� �8$���nRi�qH�->8(k�Q���M"NP@H3��za�d�U`�p`�2�{P�x�f0���]H8N��O�z���)qpt��� U<a�����"��i���p��O!g+�S� N(H��Zc?��_����9"t�SZ<����B��qL�^�,�Ь�Y3ėcY�"(l�x� ��,u�3����G��n7��b�	�r��\�� }�}�t�Bp�{��GؐLǮy�1�l�</��O2;��SA�w1������@�dl<"�>��	�ғ�Ltծ�G[0�;?Q� V��oT����p�g���>.7�S�2��E�r�����7�6��7�b�{�����C8;~@]һp�0N�&Ӛ���~�ے,�ٺC�@��� �G�a�$����@0M��T��怒m��|S=Z>��Hnɐ�h,P�":��E�u���o�^tc�~���`H�D"L޺�t;�v���IFpO'�t/9q,�bJH�3&�V�Ye�4�ʃ��({��7`�\\G����� +͉���]�s3�B�6~�غ�!�Q��ǜ���d��I��n�;棌m!>��ș����Y���K�B�;�ŗ�9/6���:��!cC��{G #���I�e��巶u���i�ʻ�x�{��ي�� զnX�x��f�D�׮��ϑ���2u�����%O�QJ<���i>b��{����y�-V���d���;��(A�%&�LQ���Ŕ�Ӄ�A�aE��)�����<�S��&�q@x��3�_bR�pb
�r��:Z՞0�cA��8�F�[#w�=z���=�&9j��P.��9?i{H�<��3����m��v'���{�o?
�hn�es�(�ٌ�-w��疩y>b�Ž�$Nꆄߪ�ُ,J��T�&�~V=�:�c��?��Ml�<M�o����K�Kd�1�B��Ư�Ԣ�S9�^)�����p|��o�iO �B���ɽ}�O�9�7��t��>TX�
�*g'�������Ђ�#����;X-�����-��&���(� ��z��+�7He���(k�j!����۸�ȞLj��j�F�'	�X����%��9�]�2���Ҫ��L���aK�vx𭠮Ƞ�bj.֭�It+;_*g�|����X�]�9~�y͎�W�2*�$�e I��n��<�>��@�A�A�,�n�_y��$��B9�d���h�5~�f��p����$\�`~&:y_>��ee{�N��ǝ$n%2�{�mY�(?�ˊ�+�^�m'LP�U�#����@E�+U@�8֪��ε��\Īu���q��E�G��R�Zxx6�s����=�(�x����=��۩�6��5:��o�L�p����l��q�x�kr$��ͳ������N�����"rs����ȿ��u��)"���1�F���Fx8e�$�O��֊�T�zF���õ��
?g�$����f��w<�'�l�q��pj�$�D�&m��*O�w3�iN'W&?-�����.����_�-�??�M��"OfI��k�n���J�7��:�\ W�y�B&���·�Q1܎���;���ub�N ��C����r��P�^�ǃ}�n\� ����v�+�Je�����r:b�Ԧ<B>��a�trA�`7B�1���.օ�c�Xч�hᰠ)��aJv�']�&������+dn9\�avGcz��w/�L��:�����0�oo�|�<����7�����`�T�.��mU���m��d�dR� I��b�'\�xY\��P��l��DuY���r>��Y�m��`�� ]u\�^����:#�ݟ�#��:vX�`Rd�cBD��f��(���Am�*\�Z�p�?����D@�I�;1E-��{���b�]I�˫'쪍�$�ݢk7"B���>����9��b��z�c�u��	�t����>�ۄ�����w3d[����$��Ш|g�`�_q��g�0j3�052D���̕|��K�d�/wOS���tfy^�W7�9�̷��C��L��`U�o�f&D4�}�ƪ�8���%_I(�]�g�#����=�4w�R�c��O�i�%9��S:���I�gE�!�˧�*���D���%5�˖' ���ʏ���Lr7JOٜ��,#���*�!�5�����;Gx��G��u'Vd�O��	��܄isl���A��Y�/c�Ι`� �-Y��JQt"����75�����(�bY�.Z��-3޾����#�Zq�dd��f~���֧����4�,5sݦ�����1�jE��v� x�c:�u��dO/ӆ0pò����$���B5�h�lN��B��Ż��L���	�呂@���D�A��|�7��+�X-��W�jt�V�!0�]]���[�f��SX|��B���6�Hʿ��a�?�S�! ��
-�Rݮ��jY�ǟ���`�	8�3;���2�,G�|+���*F�írغY�l��d/�}��S��bq`�z�yhˠ��k���Զ��k�B�B��$N��$�gh��:M��ʀ=���q���z���8�.B�T� ��B��%��i�����x��Ĺ�̌�QEԵX��K-bkڡ8�+�����IШ`�O]�Cu�E ZuL﷩9�[c���$�ῢ��f��b�z���3S!U��(�J �vA	pM�� ����a���͜�t��ݜ�U������.��pcަ4��$�m�W����V�˄�Q���5w�t�A>9Bx򎁯@k��]��s�=X�K''����������:5�Ux��Y��Jf���)ӫ�n�=E�r�_+����H �+�i������-�d�V�V���#)(y������h������K�Hm�[����aM����E74���>�4q�F�������A9.}�&��_��g�K>ȿ{�6~.F�ؘ�y�+9�^�n�S�$�Y��b���m�|E��2����[����8�A2��N;�"?���ǃg�R�\L%��t���U{�N����ǹs��D�ݣ�XȠ_�g�/4���ת?Ⱥ\#��m@W�Yf�2��c���I'�6�5~��+��Mi�7� �? W�&��S�y��f*�{\0��#�j��
����^��}
�)�oFQ���	K�6\ge1��A��P��>>��SH�o�+m�&�3�g�X�z�V1o^�NB�*T��R�fU�M��i��������N 1����6��d�������É+���-ű
�����J~�%e���*������Ұ"��	,}q	��m���8#̙ʛ�c�~c4��B�֝�z�dN�ި� ^�m�C
��Q,��x�����M2�I��q/�h
 �����ڢ�"����Cfӈ������~��c��O�o\٧�O|O�{j�tTO��`�f�6���[t��ěFPuͼKV+��ONոġ�./"� Xlc�؈�a��������,&���L��F\�Ş�^�^�2
�j@�Yhtm��p)��қ�%E�J�\�5��=?z�+Z������^ù���k�h���/��M��0�c+[d�Cu�)����G�BǤ҂���n�F��z�����<U�%��G}6^�<
G kA������P^'����vnLR��e��J��[�%�D?�e#nS���f*�I�䄁/�Ml2m~_#wJ�k��i��T�"x���~�?;X������]��^�z�����^�����^�f�kM��cd~�����#*p��	{�q���
���=�]0�!M�F�a��j���	FxEu2%��u6Yg�g��[@�d�큀��N{7c
��m�pJ6[%�)1�<ɚ�
�I�DK���O�1K�P�Q�Ջ���%��2wy��2����f2���a�0$��K�T�6�jx�6� \�3[������SK���}����X/�� �r���^�g#�?M*���Z:@�d��]rB͝V���$dr���Y�$��*T�Ӡ�������R�u�s�.^�+�,M=�4�=KT�a��9x�R����T�T$���̘�DB�L���#?��jIM�\Gy�E��H�����4Z>��mf8�-Ɇ�\>)����� 8��F���ϓ0��ࣔ\aW��'2B�T��g�=�;}e��p�JƟ�e���縋a��,�&|����o;��p�iJ�]����J���i��#���.P��IJ����	�T��_�ѭіi�VW'����߭��͜q�uR������'#x����s���;4�c�	�Q1�gq��y�*T�hC�=�A:q��= �`����Fbߎ?vS����sfR#��G������:kp�_ʡ���H"���x5�	3٫�@1���S�
]��� Y~����3����ߗ��&�,2�8����`�o��=/ґ�m����\�w�����1��_�������J(����Z�|��{=^����6~g�e?��"�k&W\�aZ���g�\�n����Ŀ���p�<����g\X���'/�E�`2�]�k{�1S,ϔ:ޅ���j�bd��BL�/j��q�LL�7��:�.X��7Ӄ@~ǫ�U3��k�]II�nML{��烓�@�9��U:�]���5�v璎��7c+���o}����c�6���k۩Ƭ�$��ע?{���mQ�:��
��:�L���p@NPzl�
��R$�!�3N�X�ɜ��L���Շ\ъ*dO	�������}�]n�Kq���~�k)��F:�ȝ�p��֔���~��ق���[|�D�&�\�Z9N�/Aƴk�.�\6@���ٿ6bǵ����g �����8����kR;eYt5� Ē�ý��e{�0�՚�� bT��Jd5=�jt^�ɘ_�濇G�� F��[�)�
�I4R�҇�|��Y�Ǝt�I����_�ct0/�]��ت��w���s��R`$���>D�ɼjG'$#M��$�:�����u�J���6g�R/�Y^	�A%�7�W��|���L���#(D���ld��`�f6(��j�ŕ0�� <NS�h��R(������(�;���@FoY֜��o��Z�tp�nDl�'A5����%D��H�q|���ݮ��NV���ù�����M�E�x�e	���$&�ư�X��3�(+C�;U�:���d.ǬW�6�4��n�8���u�G ��y$�K���Cm\�eL�'Z�%�6E�O�e�e��)�N�,Ux�����o�L�z���z�g���U�EkV@)?6<4ߔu$?��=̖9���U;/�sL���4�Q�K�j7��0:n�J�"eh�[/m�)h�)�,
�̇�N�C��4�~��b�Q!m��O!��-�H�	�[x�~��E��jo迨x��7�хjʚ�W2H��;�Nr"��a�F6˱=�,G�m�����_���he��)?b��5(�N`�Dғ?�X�����2�D�<��dF��r!�nC�7��k�"���e},xR��9S�R��Ɓ��KMe�B,y�(�5�E�8�g�)h6�9��Ǟ������oDn��&*��o��(*��.*�1��k�J��sCW����&���v�� ��W�<zM�����׺4�,���Z��W4�ǖ&/=��M���Sq�u�?Ε���%:���c}
�b'FL��|W�J�𕫚8�u�vO�m����"��B�>��'�=�JJ'���d;����j��Wma2�pPꀞ�^
O�u�	ϖ�v.
��D��h���3h�͡����j�5�N���)㉅@�~�Ȟ�eW��.���!�('�)�ۍ�<~�r���D��9U_{m-)Бq`l|w��l[뛂�>$::�+Ϻ�1��&w_�-�h��C��:���Ӯ������%z��Fh� �єL�e_�eeYqS_��fO�8Rw��@)v!ZA�96�WMUkb���\	��D�j�͇��^̟��ub��6��(�Qȯ�v6,��4OE�YP<^��:6[(����k>I>��򠯱^�C�Oo�ߔw�u&b��~�؈�J�C���>�`�i��-_��7^W��K8�]FR<u�׌���InTEO����Fd#A�x�^c��-,�ob��-�R���N��"��5�VAo����/��U��լw��n��UY���&��A�CpW��7���JE��-ͦ�0#�-}޾D"����ձ��_�"d�@0ɧ�FXT֐�3BR!�g��N��4����<"tw�N�\l؜�csn[q2�Z��
���+���VA�4�
��t&≲[/^=U��K�E�f��CX)�ե�%��IH	x��Y]�Y�8�+�=Q��(4 .���"R�-�ɀ��^��7�I������Rj���X�9mzEL�"*e��/g�9!�U�O�x��G�V� ݑ�\\�f r���0���Rs�8�b��e��K���]���̟JQ<�W��n�;���/n�݉��
����P��I�¿�����s�1Q����2�{���n�ֶ;���o�K�
A�ǻ���.��pڙ_V����Φb%�퍚�����³���7�����qB�m$p��%I͡D�"L��^fٙ��W�[��J[�=C���"5�.��#�˂6mS�� �46�1T�Pz=Ӽ�n�/s΁��jKS�P��Co4uɩ:�0'{N�e�-S�>�V\"��\�7(�j!�Ϋ)DW� ��Z?�vg5�B.�b��CHW��$�`[j٨�,#>q������јYt�a������kH�� }�Q��	��r^�PJ���{f缁�<(�K�B����:<,�t����Pl���e��|��J7�����	sz>� R]����z��wi�a`�;�U#�>◡��U��`�������b�!�������I��4�9^�:I�ь6���5.�Y����OD�Y�͢זP)��(��Z��	��I�W<�۩a,F'�\�t[��j��rb'�T8A�ꋂi�[��fHW[���T�M����o����	�B������$��,��)�z�8�$A%�G�������K&3{�i�H_��PgJ;6�e(�r/���~��d�u���:������[��|fͼj�G���7�����,�W���_���k���%�ɤ�;�hwx0W�!�L.�(O;�����<~L���@Yn�a���y����O7��Xc�͆�&T����*��x�T�y�/���0-�[5�]��P�P.��5l>(v���"��x����~qY&����Y�a̓1[08�̴aj�3T%�\I��~Q'f��]w�}�`���sE�&_g�P�04���K�L$��Z-�s��L���&(s���y�慲,5~uI =a�Tg@c��)v֫+�^�I��ε��ќ�<'C�g4��E��`�W����*�-��s&�v8� �Y�����J���E�̀�H7ɲ��۱���fB]��ʪ0�Y��0qM]�*�?��/�R9!B��!�����v���ym�R1�ǜ^"�Wy�*�}�ˏ��j�Z�c��v���po�,8P��0�,ϔ�="��P6���Dl�Pd�Ř����m<O3
�
�p��K:�i��!ϰ�� c ���+���$����<�f~�l(����*{GZ�����§�p�ԉ4��nǎ��-W�������<�?�	u��N� ��ɹ����O�4��`�+��V+����&#t3�z~��Fq���k���{����'���L4w5�^���R0��Н�1�&��Zk��ֆ�e=�>��d %�A�!-B�)H3�vTtW!�
B:�L�)��S~YEr����+F��A��Wv�� >�!��>3,�NɁ��/&E`' �|D�v���1�[����T�2'��Ir1� )r>������8��$,w�yc���q� �*|3�>�Z]݌��Άz�u7�����^7��3s�-�0u�k�[��漜��B/�'K��0�>@#�́��M煾i�ġ�l�z�a�]V�J-S�(2�ֽ2�LKP�9�%z>����p��D �q@k�-�%�GbA^*C����gUk�������4%`�N�x.�%�3*����}��p߃B%�;
#�C#�?����Cn!�N��
-��A^i*���)B{�'�r�B�s�>����Y�{[촢��<k:ŕ-�þkea�.��� o�#�=���ԒO��e��l�\���<��J�o�;�Vo�;��Z�g�6�E�mE�����W2�}�5�?M��꺎K3�M�����0wP�.����rr��U��{�7�;��e-���սE2l-Hi���BR9�"�ܜOf�ܢT��OS��´6w$IB �%���<�{�����h�i�Aw.ɔ�	��K�����t.�*ٚ�+R�s�X�������Fűq��/�2|�mQlt.��I��v��~_fe0��S�Έ�6�]�H�����
? ���X��F�g�'�m2�Q��h!�5X9����Q�ҏEЀ�� �%x	թY�*D}����9�AC��ԡQ!嗩��,e$��1U�8^ۻ�vu۰ 4������ #;2Q�
�ŋ���C:��L�=T{ʧü,ByRœ���YM�j7�\��F�_���]-��^����1�F�Me���#V�'��_�5����#y#<�7��۳�赗��@ǥ�� �7�1��qᱽ4鼘q7����@�h��\�hݲ����q�lM �%,�!l���+a!�fW��FՋ4�gvy� �7��X.-|�����A�)�n*Yf�[���]���2@^���N��z����������H�Z��r�`�A�̺����d��TrF�ӵ$��=Ka?4���9i?AQ����A�c�]WS��3_���Ὧz��LO�{��]�D^��ηh�u�u:�R3q��/�3�����ћ��J�2����#���+�y�	luZ~�JJ�)�@L��:���y��JkQ�H�-犐p)k���9���bh�|�/T���Hr�CYVe���Yk�|�݀p
�!���-n>�f/��ok쪇��7�[�
��7�Ӑq�VV:�����9ۯ�����bP��!zwLZ��	`@U�]҃=�:f���<��O1�'����PzP�xeG�@����䑥L�r���W:]E게�vXϣ�_,�� E�v�	jA�Р���֫D��5��<�u� 8�}-q��te�a�處�nF���\�_��hg��|�6�m?�ôt����+~��������o����@���ڧ�"(��>��E)��Ȑ��	L�t���/"3��KecK&5��ͺ�(z�N�V�l�ˆ�V�Â9��ѐ�/�f���T���9̿��Ȝ�W��-�qj�D�H�U%Ih��7��p�����,��4�\�h��{�!Nur� ߣ�|W��������P��ذA��!���1pa>wG'q�X���ya�'�å��Fr�HDw8�mD�ƱY�Rq�}��b^u�& %{ F8�BLT.ɿt����pB�A�_c=���}�#���y�zd���0�N��H�	�&�{7\�*I�znG�8pYq2ң ���)"�f�_��"wT+����xdc:��~�|�M�֕>(7aj�����(�.V�b vPh�;��Z��6&�� (O����a9���쪟��Ρ�#0�އ���f������_�۱r:{�I��gj�]�`�w�7!��C�܄k�<i�{�(CE�ͫ�� co)�?˛�jB:���`�MD���c�#�t2� A��������w�"Tt������z1?ws��ỵ���#�^T�h�eNfn�"��漝?�.Në�%H;B�vr5|���Y���҂�����}�]s-���8�{��ɛ��b���
�'�4w�׆9'CIS�}�;�43z{��^��R]�j�B��}N��t	� ��սK
�^NL?�9-�5}FV�����/�e/�j���s���i;bR��!JK�1��:N�_�m�5�����u���#;�ed��u�+�V
��q����kf9k��y{�k2���zS�t�gJ����f����"���oű��J��(�"��D.|��y+�������)\�����X��Q9�)�/�P2E0���� ���ؖ���i��:R����U�ڣ�^��iߎ�7�^��`n^s��#U~:H�h��M�����P�\���"Y.Q�=p��613���{�����i!S��}!8H���ޒ�\�/�-���TZ@�'l(��q��@���<	���}�~�ldb{޽�~���l���;��<5d"�1�������?������Nnro ?�ـ��4���{zm�g�0)}��Vpl4B�.����L�9��feۈT���4)+J�[-H<�b^�z�K|t�c!��R�HS�Q6u��L�4D$�t�R
/ͼ�̯Z|�	�ꉟO�#U��������&��~H|�K�L�yq3��H\�8�+2�`���n~��5���-Pƽ�]���<&sH���@�t��K�$Ë��n����;���U�X6Z�:�Yk��|'t�8.���:I�3�Nnp�/=g��i�vH	�6�8����Z��AF�I���J�p�%�4�ٷ	����
�����m��f�0Р!�����{�9YkI�����̠��,D��P�;)��	�&�����G㽬��O\�-�u�.��D1l:*,
�'g������)G��1:}�~U1iI�}$8r� �8�8Z�����z�l�d�T��Ė��Ou���$Cƫ��o;�*_0K��%� ���T�v�E> ��u�k������P�q*TD��p�K������ŷ��r~h�)�����aw�����,V}{�k�D�~�n�I4/�Hh�S8KW@�d���.=2P�O�p��;	vpSo�Ε	���T�x��z�A?ʱq$��SE��k8s�����ʰ޺"�rϫReX|U��}��k�~ҴQ�z�OɬCd�%�p�VO,Y������^AƎ��2�~��xԌ���
�^UI�ۜ�FSа�u��vŚ_5��F�X��982a8S$����w�vDa�>��������i�ê}���:�G���6"w�V�;�`n
]IH��<�\׸q^n�y]���З�@�p����h�Z��}�=��QHWyM�N�!���UEh�1�Bt �97=F���07ù�RnZ��·mǝ:��n-�?�X�Z��0`k�q�!7��T��]�a�Ŧ�L:;��i�9��j�4��def���cj���r.N�q��� �3��R�f�~�O{q�{0��j���w��7�~�u �I��@H����A�x�}6q-�l2ǣ���~+�p��l�����+�6[�	��H�o��� �s��C���>!���8h�|(��C��{��G�A�:ّ⌀\�۟A��f�d�QBVy"4qغ���/����0�y#aԥv���|O�`_�>�}�(ݿh]��������/P��������$�V�o];�6���쥒���я9���W{\�ԫ����39j���;����	�Eb��&${D7��ǋ-��ޯt\Ԝ��k��))���vp�p�t�O��&^�������^.���qkA{i�@��g�9Hg4_�:|�9qՅY-���m����(��l�?!z�R):LW�y�?�%>�o|��?��w�(lo"A��u���F�@aN$ؠJ�"FRp�{ @�u-�����1[U�Z����Eh�z�کXOf��{gɓ��L�3QP��
X�.�UE3�&L�x�Df�ݿ�I��g��R���Hk�����B�
�_'�ye'�v�ܮ��~�3Q�+��Z�^�@���U:�D`���6&���.Jx#E�[��&pƐPa6.m��Ѡ���~�h�s@4p`��!����ԯ*utpZA#>��V�����RԪ��\)�I*�sQ_�G��s髆.m�ӹ�`��݄j���A<3!���J�c���y࡯���v�ceul��~��(���������h(#)a�L@W��<���f�#��o��h�\���qȨ��Uy�{��.��|�vl�*ۇ���ȁ��V�z�$>W�P�Ǯ�jWY� ��ad�����CK�iC�e82lb��#�Ϲ�A��n"͚iH@2�;�:�{=���P_G�Ȧ�+�P��@J�)ţ�<$��H}��G��ƴ��,jߙ2 o;�"�#'qAg���v4���Ga�����;O�p�K
NH�?cz�9@���c�'��7�ӫ�R�������#3j�M-�2s����MÉ�a%���DJ=�<�r�F� paSl�Օ�5� ��?=rS;,(����f�� �e��ԹM/xx7Z�����9��bK�4Z��>��n��	Z�`5��wv
{�T��W�/p��tYd)9L:T8bH(��?c�Y <�[ν���z�6�`��f�r���9��������աe�y2�d��V1�'5�O�ף��Fy/bq�J�B�� 9l$L��1��������IE�����@��K}@�ҋĉ���/�h��#��T�~/�s���%7�!ѪRy��6,�����S�ξ�Pޱb5ös��Q���
�!zQ���d>\R����k8��m�v}�qF��:d,<�-i x6����΁�H%x�S�c�7���:����}B�2(hY�6"k�7���ge�/�A��M��S� �5����#�h�Ҙ�|�#Vk.Sp2�x-�=��%@�M�%7���n�1����g���z��tI��I���������#�.' i=v�6��8y��|�`�j�� p0Jύ�D��#np�t&���LT7@A�n�-�����G�;� 	l$��0�ˋ��(J�˺I����y��뽥P��H�QQ	YB}�"�A�; 9Oc%��s`�c��w)�q�&�}�K`*��?rTy���8W��x��R�jR����%��HS	1C��|)�	K��K�W��cפ��5�X3l.�~H�AF[��?�w,�/�_e R�Q늤�LC��%R�_l6=Q�!��'a���P*c}>�q�������vmp�o5�ʹ�z�DFTgE�^����ư�j]�_Crh���!A�WZ+�#�GиS$�sE�f�+ޱ0�E�������V���^�����_���{��#�C��<R$
 �,7ApO�N�v��	�s0�$`tv*=���Ƥ�ߛ6Z�({¼��8{�ޣ�/�h��x��(ͽ��SB�.���vE�¥<	N�������� 馯�!���u:P�el�S�l��Hp����S�8����tl���<̦g�\(rrJ�u�_o��]�E�5�}��Wh�Q��F63�,���]ѯue��c _V/���ɬ�?�>�)6�7/�4�Pg������
Yv0�R+��*%���|�9E9]t&A��)q]I�?�Gx[�����j+&�'I�9�������:!�d1{��b�=�_�f�3�.�X妞�n�C���ŏ��+WX��+5��lEq�C=�/��Z��ޗ����fn�ָD΋A�� ƃǐ�	D���o�oۑ�&&��t ïA���Nne,�dB���Ř`�
����j㥜mE�͍,Qmt�slx�)����K�8����"�~>��e%V*�[�ŦlA|�����F��˽��$�����^��'@<b���G+Q��;5Ρ-�;��"%�)F'-��^�0��`�g/�>�c����j�;,� %�E��ɂ�l$(Թz�W��*V5C|���@y�ݹaY�7.�y��_��]�����}2#����v�Ͳ�,pXY�����ɡ�\[��xq!�Ǵ~��%���B�{ {/�/��rߞs��w�yH�նF��x��֎Z�5����g��5�l�#}�:xkSV��\H�+#!So�B}��e�;}�T:Umg$ㇻ׷F��^��������)a�/Z�!jH~�嬓�<�Vz�
���g�P/!Xk׺5��4��/d�59
@n�2�gc+y��R��ڳ���nh��"��h�$�yk+_"�of�)��tΜ�[�qo`^: �lǺ��)�Ca4��W:�o�Q�둛�Z6�l)��g?�~��ES��,{@��Sˉ|�7b@
w�"T��lF"*�����Rn�[��C�)��*�FŎ��o��Й^^dcD�뒙>:w7��~3�-<�D*+�����2�3�h6��n�++1x&(���C�%��-��Y�%���ߌ��?*�X�[�a(�!F�6R��L&7�i߀;J��n�F|hm�3Y�E�6�ęKB�;����_88~�)mAIE�F�D�sj�l!(?��<ء(���$���&���<D|��^x�BNDם&�ȼj��,��vr^|�.��q#�7�-Q���hŊ{4�����k���"�ge�i�q2@��q�Dr>8<+ߕ���i���b���S��2��vg�V���A�XS<��v����Ge��m�p �Dh��(�+�C3	��g��}Gfve����$�6A�������'�>�����2��ts�<h�O��N�V���e=�j�]l[pZ�U7��M7����[[�h�b��a������ү��o��X �e��R϶]�>e��8Tu������
/. ��f��r�e�@p.�@~7�ؖ�,���� �# �d�
�G���c�"�<k;C�P!%�&3���H$��8����w� ^���0�|��Ǡ-~ E�Iݒa��X��+Wg�R��W.1�^�Z�xPg%�"L,�7~�
���sc�-.�zI�M��8��M,�qXsA�kI�c�D�@����	�@R\d/��uk,��Rlz�o���L2�Չ��`���ԏ0������wNP��Q9 �9��.�\e{Gg���̴1�,��sNԕ!Q"p~��$8Ԑ�G�;Vhb���o���'�Y&B����P蹇p�k�����X�|G���u�=�������!���"�T���m�ߌG����UvEBO8=�n3���J=pߕ��C��$�S��Qi-����۝W�)��ʭ�n�Oq���7�����0�e[��}�Dğ��L�PUS53���:=�����&�BG#����?S��w��_= p
��Y�^)
�jzl�,!^<-�4f����
S^9��2�5�B�ʜ1�;�W���¦��
�F�D���V�B�T[e�~s����,s��G�"��B}�w�=�@--m��\�*��djR?;���n�4���=��?�Χ�ٟI�ĉ�}�k���M�/+��)�A�)1�,�E��z����^���1u����ܔ�ƈ��d�l6Xk���I5���}D_Lǳ�7Q�}tq�ٔ�&��Q�S�y9��/@��H��r�N�A���U� &���1�|Î4�lH�����ѣ�.
�K���d�Z/��C�k�DES�S~�����b��j����%���wf�N/�rq���=r;]>~Fǔ�,Vp����u0�54�U�v��S����P+��%���n+��`��C��0U�D��_C��2J����x�	v��!+䔤T��eIZ;]�h�p���h�1V$o�8gW��67��C��1pP�y�C۰iͤ�Fbg��M�q8f����m�gK ��E.�E����ԲJ�� (�J���g��P%�ﮡ4#���������D��	W�
��0�[�9�f:T������c�8���Y,n�#���ۇb<`s��$'�=� P����	Oo�a����c6RG�hْ��c���4'KL�zvY֩qi�)��6��ĭo[�1�Z0�ZX�)OO��\o�+���b8���Ŷ��v/�?�d�m��۹Q>�L Z��Gc�X�ѭ �V��*��׵DG���(Y����r���u=������O�4i2o��#������[
�Wq7��G��"��*h�Q�]�����f��:���;��U��y)�K�jD�g@�������8}	�#�{�BJ?e�O��WX���l���y�v�u�/�BC�ڹ�9S�����	����BKxE���M�v��V��/D��keP�<{�SO�LO�p類͡>���"��yCq��ؾN�NI��i7���@�$qx#	ݛ�R� A���`��ء�ޫ�I����OA��f���������%@�5���!�5�
A��w�XzY٭I���S$ˮň���)���1��-�_�C����sQ�>�ׇŎ���y�-0?'п9�5[	"�Pڗ�J��l���%�=>j:�92��0�F��J���N�̢޶!,_���O���!��w�łպ��ğ�:)��ř/�o��q�ϳ��M��ĉ���bɽp��0���К4 ���^T�e1�&,)X�O|�XS0�L�E�]�DV0�G
�h��w$�ۻ��$�������	N�(u
>|�R��wx�$3i�1�V�X���������j,�)�#Y?���@܆����Xj��Q'�-��8N�9/jKNL�0q]�6UE�Y�X�'-�M I�4����� �I|���}�N�g���H��S�]4�0�@(�����	�	�����V�\̯R�]X������:�N�=:�*�D}iiK{|�^��e���q�O���CO� [a���y��|m}�m�O���}PP׭
��=��҂�U��uR)ںAS`��k��(KY��t����|���诏���I��_pC����)m*�E��x�PRV�s�~6��Y�E�Z���B"vtL>?ɵ�m�yE�c+��w��'~j�!@9��o�Nj�\|�[[A �R������(����ǂ`�d�1p_�E�]q�K��>d��N�Pw���@;w�$B��s�Ѐq uh�4B����_G� ��:F4���t��,'��NAZ�sm�c����j,�j�o��#s��wH�O �d�G�q�S�Y�ؙ'���s�eY:�}!w6&vH-�9��i{�$�)�*	��^��L'V@qʤS�y�����h����P\D3�B�i<rg y'����R{�ƧK��61����&�z�p��Ho��ye'�4��P��G���Γ���l{#_[���a�&~�WaHs�d�ID���;�Jٙ��d���
�M�r��Պ���n�`Ӟ\�9͢�;)Z^�RC$�p�O��r�"�&	���,�2?
��q\O��山�k�p�P�et����w�?��Ћͬ4D$���ן_Y���^w�� S�����)4);���&�ư�+��[��%.T� �4�3�-�u*���7�u`N����,E�Q~�*�3`*;G�u��Q�a#����]p�v��5��%Z�R���Ւ άL/�F(<d�3�mI�a��azΏ��t�ǻ����P�s��ϑDb=�Z.7%�J?R3�ݩ�� �<�<�(,Е������]�ɥM(� $G��E�ü]ۥ����]�lOh枒r��D`[Pt�
 h�`jхl�������n�3�>�@s�K<QK�
�M���Ԁ�xɗ>�� �
X����G P��?F��\٬|�����L$�G��&����E���MT�g)h{̖�o�����Us��v���)��~���v�[<�ϻJ�4�SXQ�v�8¯��1�r�hou�n��x��
$�h�\|���)�br
� ����p��|����\���@�����}�^���ul�7,ֵd���e����%"��Jƅ^�,[�#q�Q�
оA�&Qc*����Qt�����腆=�}x'�+Z\Y"����!�ќ&��������H�_.�v��(�=[��YJ��:~!�(�)M�cz��8p��|T�������t��P.�q�7ء$�䖃���b�AJ ���Ǌ��|���
�&~�ȻO�J�b���"�/� dsy��BAQvs���q�.
5;�v���v�(��ٍ�S�,F֪�@�=��tc0;�����+����}G� �*m��c-0�DάA��^���j�����:��:�/�����4�jT��a���B\XnK^v�4;ծ�W�S�m���[~�>|kTJ�** F�� �IZ���z7F��£I}�H\��a)s���&Ylkt����ھ��d�b\��!�"R{���D�aKB�	8;d�Nf3x�6?�e�>�a����u�~'n�6%%m䛺��ɉ�4�y�d�M�a�*��rW�@���C%ZUCԣ�U����8�r#�qR��`cl(JK��aؤo�p�9t$�~���p�&X���>�0��h��uMd��8�ˈ��K�G@B(�va�#]����3[8/�H����T�8�Qk/�r��ݴnp��l�:'���
p۪���Kq>X] ^(6��2�_�&M�?�Y2l�o�-�3���ׅLi����2�˭��J�ϭ����;g��î�L�J� A(*j4#�Ե�69<��ͫp�������t����M+װ2L����2�H��B0n��NY�J������8�kܫa��*c�֌�]%�����������u�������O`�P�S�{?���d:$����2�}cZ�K��{uS����T��!H�U�K֞V>��-��R{���m	蘊��ޏn�VJ������f}��.����'���ni�(��'`��gl��E?&B�qe�����|e����_'&��wNX��P�9 0�R���)����<'!
��Z_�j|@L�da?�1YhrT�����ho[�W�M4']��3k�mDQ�&�x�FH��e�����fQ������q��.���\M�tf�ǒGv��#�İ�ʳ{/�8����\z]+M�
��tLU�.�?ԭmůT�p��\�-Q���8���
!�f���Q�sp�Go#�پhe<�,�ïӰ��d��
�Y�WD\[�)1k-yf���%�`[�rr�C�-��� ঠ�c��[��� P$Jb1���r�S<�6���v��U�G~v�ɣ�H�����#�����A����@����(�Ȏ�z�:&.K�6V���~H�VV6D��/�]p%��C��d��{�}��ȶ�
խ1�8�9�;b$s�P�M����'Y�we�غeI0����/�U��\���" ��@ �A�p/`��-�)X�e��A�����+Z�L�ŭ����&1�����?�缑I�ڕ�1¤��%� S/_��Fa�ٹM������>�j��\�̛�F�b7���b�桶
�9a�o�#�h�}�:eGuT��C���h�u���]�d
�$��j�׌�7��n��%�f)�,�cx�[B"ߍ�j�^3LlV;2ADb���"�w�g�]���m�F�*W��b��2g;Q+j\�Y!��V���������:�Q���u��\�Ѣ���OZ3�C���ﰺr��f��͇���M�4.����!�L*�]�=4�Ng#� �Ð��97�;�)ĝ 2>�;Eq%��b�b\��W�v/���s����-e���?q��C������KQ	 �9��xj����U�����& �A�R�my��<�����"��ܹ���PJZn*l7�J�t䐴F%�|��NqU��=�=gF�v.��c��_�F��(q��F�b�v��V�� jL��BKnS��O��[�N� � �ތ<��b�2yƎ��6�uo����~5��-IC��o��cג��+�O��h��6=�D��=4����
�Je|M����o���5]�����r(�A�f��.-ҡ���d�v*��+�E�W
��䢛�b���wj([7�Mp���P<8���8��Cq#�v�猌H���|s�X>V?�6r�[�U?�>ѸN#T/J=�^'���G����n�>U6��/��o`�6OG���p�6ym�Mf7���W*7���z_�]�~.hD�d�[RgJ5\��� dǘ)3u� ����φ�M���m��3R%*dh6U7m��ij��/�D�,���8m� \���u��;�Ih����Z0�c��j�,�=.�)!�)@���LYѴ8<���SN��<E��MSv��������ͯ_vc���<��������
t7S����;-#M���ͺ��#&ctW�����҂eǬRXȘʱ����17�Qk���kJ"h|Ez^Cf#S�C���M�9D���]�ߙ5�<���Ǫc-=IwD�Cl�~�5���;5��	x� �o�͆ܠ��f�&ޟ�|��6m�arR ���^P�J;�y��w����8����RG��1w��B���"��^12�����-�� ���Il+���)�Z�Q�{?Z�i��&9v]*�&�^����L
���:�z����ϕ����k�|em���|F 1�k��K����o4�`3v�6�n�?�X��@��j�˜�~
�Jw,���}�|�� ��\�}�zN���q�|����g��qx�������4�P�lq�d��:�ʣ
;�K;@n��Т11��J�m�Q �t!a�?oq�<�o7���օK̽ap_�`�{hx�R}:�Ǐ�r�tm#�]�*��j�����r�v���< 8YN�^,�U����覭���񸢲h�M��yi;��d���j�{Do��q�*��3o���K�/$�{�����y�U�;X%����p6�B	����
J��9�*G������ۻ��<['���R6���ۛͯZ�hG$���u헳ح�R:O%_*	U�Q�N��FY�;��'�~ƕ�9_d۾ъ�Ժ��O��{u�J��r�V�$�Et�0!�D<THhI��]�p���%guz��*`�Qr,0�ZE��T<��o�w���3R���K;��K���2Z	�dp����(���Up�5ѩ�,w4�՗�>�,6I;N�jR�}����aŋb�D{"��p�����J�b�fxu6�5�d�����9+�Oy�P����@���oQ�S(%j��Eba�U�Ix_ׇ�G���|��8���B鮜������2ͷ�#��]�f^�n����kn|�\Ȅ�6��s	ulU�B:��xʋ�xG�pM)��s]���ԏ��1�*A�٬z	a��̃t*C(|_?4��|�<A��lP$��	��m���^Jz�%�_��9/Ѱ_��5.<�� m;t.�"�s�c~��o�����[�f���
C�I�A���<ۣ_Ig�zr�=�l�>.M3M����AP��t��P?��%8Er7��M�U5nk��GF�*�e������Tbw����?�:�j�c��0"�p�aϟ�kYѽ٣����6�J7{���]��\}��6JǠ�5nj��n��߁�2��!0)�VϨ�h�s��.s*�2*H��T�r wz$�E(��#H��r���T=NY��@@���k <���5�bB��RP@�s�qx��"��u����z�a!�L���0�����'�Z�oFg�f��m=�bFO+D] ^���N���2��-�a��kװg��f0@��;еv�	���:uW�6/��k�4��<gqf-R�R,s`C�� 1����ҙk�ɕ��C'â����=� ��Ie +�#�J5]�T��J�3$D���C\ō�|�M��j����t��9˴�R�K-]<�iq��s���eQo ���I��u�}�����]"��4�ۡ�!��'��\���.���~�7{A�I�r3Ϟ��$W��m�D��E�Sd��Q�c��;��ɷ��E�w4�<{�[Z��p��{(���A��zQ��[?�iG��dP�	
�?�(c��N?\�ԫ��Wz���R�h���EH��0fd�����3~�LqL�ĺ&%�o�]�UQ#�3�;�Sт�=X��"*Ǣ	�_=�S|&M��hQ�h#�.��,����%����h͉C�߲�����d���f�z;�4@�fX�reٵF	�6u=���ߦ����B"E�.s���|
SjOJ/K�̿:���a�u]������x.�!�#�]m�9�=۬����Z�ǋ:;D~�2;_�4⹃s����� 3յh������\tfM@	�/v�^o)�d5 ���8�j�,̭�,��b��~�HKk��P0>�"�a���Q]eR��7��UY��-T��Pv�����u��,l�;=�� �>=���/Ɯ�1�|X=��lv9�!�1��������Y��'����ٛ�d}��U�k,!9p/k+��o���Ǻc��������?|l��8lǯ�6�N���� L���nB�X|̺�P���w�T]��u;���6Ӗ�x���Tq_��1f���ĞhۏJ
i1R��r��[����׽�	 �j䴢����ǅ�vc.Ӝm�X$$2F��'� t� am�����w��lU�4z4F�G,�G��oq�Sq]!�E��ņ �]}�n��Z��@������)t9D5ϸXp
�֪]>�^�jF�.��A�z{7Mpɺ�S>��L"cT�'եk������I�q5t��\D�G�^]��c��w+*��$Y1f%t��=ٺ�dw0ݼ�i�i���:4�ૌ���yx�[
	����TyX?I����nf��3�O
t�X>���U�P��^����PMЪ���3��b��ZS9���,�0�T��q�d���&'u�lB���rQ�R�qѭ���c���e/`����YP\��C0z��O��Dz�&�g��;��Ƿ�_��[�f}ߟJ�����A�g?>Ho#D�'?	�,���Z�IH�k*�X@G�����Q��?�?E��0�-nc�)=��P�WZiYU'Ш��ㆢ��^�'K��rphX?)��W"]��2\���r3��J�!���
K69Z継�{�PY�h?b��CB�p\!"�;���	�	����w�u���~�
� t��\�M8�:gQ#��{:���0\�C�����菇���W���O���£pUT�����gw��E|'��.���v�;�.3E�f�++xn��~j��զ2z:�}
 ����k��JG1��략-K;P!��P��T��C�c/��%w*Sa�|�0�ڹb{�3�T�+��`N�2����A���غ
^�@���?q�ְ�"�<7�����k	.:���t�:���	���_�$䭼lW��'#
̸WU+s�D���/ss;�Fōs����]�kM�_/ɇ�����G��`��6��-��&AQ04ʦ�WZ�sq
,�n%о{:I� EUySx�
���_kM���C�Mj�1������~6�J�_��V��a��#�զ���<t�!�#rْ��"\$
�k�6r ���aO|
ݖ��&W�& �y����2�X�Ͽ��N߀�@v�7NQA/L\��ڷ�Q���>�l
�c�!1?�H�
�x�ݵO $�,Uc�?���]k`�s��m��3Ur�}���|J[&��n^�]��-��	����|���CM���)��i�j�<S5AR`Z�Y� @�AwD��	Ts�9� ���h~�䶞 dEmj6�a�w`�x�O�`&���X�q�i]*�{:oq���ȷ���h��F�\��d*��ϝ�zI�;p�7������~=ܵdtr��\���o���\�cy���L�Ty4
d_��z��^��-T����&� �ȼ��WNT�|���#�D/�r�GF{n�fަ��g��hL0���q�[9��2V\�D5�=�q.,u���Cn�~�FU/��)���U�4j  u�R�0q@�b�d������﬑I6�J>��\J���<��hΘ��Wc#�Q��b��it�z�~�ͩ/�X�`��_X5-�������V��֮�7_4'�z %�����}���]�w�
�f��7��gjs5���x=�_�������>t��UuLr��|
y3�$ [3��UHH�;ݗP�Cw��R�ob���)�h./�uE5ɶ��)1�3���IL��8��<#����ί��n]ȇ�={�}��*4� T�r9 ���V{iS�'�+v8N� �[�N�� #��^P����f��:+6�9�H�Wr��[TSG��u[�,��vr��<3����w�mNOΊ�c�/M���!���A}�xҎ�>I��|�C]£��I0~9Iÿ�Y^q4&�L=��C4�eEܪ2~��A�S��xV�i�8j<0�7�Y��z�*+�売�og���h�
>��o���O�� �=[���X;�C��uO�"v�� a1HGM�'��Jlެ���tZ�����vj�F�[�\O1�1Q�	�Y�����-0$�s8���������|�o���4z�6A{Cߤ���7W�����zꅋ|��B����z����/�v�?���A�!���Ҩ3���I�]���R�� ޿��5���!{�o����В�[8�5�į�F0�/��2`8.����@L�v��	ͮa���2~���q%�a0�4�D�ۈun j�,<*JJ3�_���jD=߿��0��2��X�(!B���X��Na-��+u~�'�-Sh(2�q��2!o�'�TR�Vؑ�1T$J��>9"�2,�G{���$��x�������A���?� @�R�l�\����6ϟsl��*�D�ƃ��}mpMg!�ēPؕ-lgr��LDF��fD�5@��+�v�u>���6v�S�� :��.uQ��y���KE�l\�)Y}��S2q��53�YنT���扗�ۥ��I(�{F���6LRZ�t:FN�0[|w$��!x�>#�&i����$?5��'d��.����W�IP|}>�B�Q�>!�$�����$��
��UY���q�U��N譎���g ��F�1ul���܎�FᴅH�Ӥ;��d������Ah��3V��3tOM��{6�6m����h�Bj/ŷ��������޲m�70~a`���J
������ݏN˥Иq6qgm_n���i�*�㕫 ��J�	5I��mWl�ix���B1�cI����3�t<z~���^O�,ی|]�P+6�5�t����������[q�O&��I��"�Tg �v�4H�d��mRNX�+���h�#r�"��E4Y��)w�NI,7{�i�}����ۭ8[<�J�hA4Q�D��B�.)�%�#�Ac>,!iͷ7-;z�����4ۍ�#ͣ��Zw8�&��tz��x~�X�[V�_Rm�o���ĪS���I�Ԧ��.�G:�^������
:��������}��'�k�^��s
���-�K����
�#�Ou�?Ӓ��*�Q����k�H��B�Eل��f�fJ8sd��J��h��WJKѪ�O�%Ɵ��~	P-��t�����^#�瘪����3,���~���ıs�Ά?dOF�-��-����������{D7^cm�_LT� |!"hέp;����oJ���=�l0�7m/�mO��>8�9In�
��m������6H��xj��Z�LJQ
�V��# �NA��s%�OҜ�o�|C��R�#�'�����{�Gw����Fb�_��
�X���2����I���Л	�z+�upv�sy��Za3��P��]H����*�Y@VW)�n�6Q�V��:�Ky���)N����̬ ~�E��!nnrlf�i)Q`�����N�D��ƆC>��j�9��m��1 _�f�b���\F@�q��$�Hh�BR�����߭��E�i���+��wMF��~���D��DT���e�?��b�&dY���K��\�X=�o4@S����!� ���}��r�NX-]�Cw���NҴ��w�����|���_�We���%�ڈ��՟��|���"�L�J����W�U!�Rc �-ڊ\�؁�"ן��tM�&ӟ�}k��9�6�n��~/��%	����B;���̴�YFhBu�,3cMy���h=&p�Ol�Т�><���\ť&�;:q��\�v��F�n��բ4��x���b�:�_�s�w���	̈;KZ�u���Y����S�%P�~";�����<�M��f>,��'9�����+� ��ӝ0�7/w�y��F ��{`�<�ڽ{�H��(?9uE됄��AQ��<���Ś�$�窯�}c���x���շ/�Z��V}�3�4s�tT�+v�����i�$|�"�̅�n?u�n|H�3�
�Jc-w��o��/X�g��K���0�^\+B��m�����d�VY${�������/g&�9��%�n�ԶB9_��c�aGf�x��~�rv��_��;&/���Tk����g�,tr�,�k��Sw�� AZ�{��YcDC|�hW1_鍝�rԲO�Ӓ"0E^㑨B�r��6a���F���>ᬺ���u+�c�Ŭ;hj�����9'\�u���p�Sg�SK�ȫq	v|���V2f�{z����(w{�*���$���B�f�p�&E�����GoLF˥k �
��f�*̵�,�ͦ�u!5|��N��`2���W�3��Hދ�]���n9A���v�9�t�=5
�C;g�%��R�ٗ�8[~6���N ų>��y��CF4V/�Eo�(mA���B�/�(�{�خ�g��"����"�[���'�m��! �l��Q1e��fЦ6R֫����6wi�^���5g�Vz�'dփ^;eP7/G(�r�
�3��ȇND����U|ص�;P쮣ɸ����p{���.^�jH�;d��Ulk��g��3O�O���\Y0��o*�1����ù�@J�%y�¦sh��6��U�M��c��CW��5eY�x*c�Zj��/0�[�j{�9�����k�U��ғÿ;��D�kP��t��t��Т;�6Z4�q�8>8�%����T@V�>������,^|�,G��7�����iiw"y+谹%���M����E*�Q&۱3�(�J q:��Y����w��Q��i�[ƞ�]��ucv�k��j�B�R���|f�#u�$���&�.h$\1�U�i=���C���B���I�0!�G�9��iv�[Z�!%!�c�?�\�w�Ļj����.%p��x������=l��MEr^�jg�q�c�I���͵73�䀏<�(��Ƃ��{Q�ma�j�'��Cl�dzp[������[�	JyJ�v3e#Qh�.��ǔ��� ��*�ɡ����2��`Om��L^��n�spdk��X⅕�g��{ ���y��yJZ��O��&CѾiy��z�D��z�@�C2%1����)c�D�r��'6n��?w���T�L��Y*�����o��0ĺ�8�AB�����He8����uDn���t���;�x�߄�LX�1���6{O*@�`�ǥ�AE���X�I�<5eY�wߔTث�IA��?pwV�-��N]Z-��dkw)����po�� �����U�l��g���	�$���3��6l_��t�dq��:���d�W��d��T<?��f�P�i��.�B����8H�
p�+SL�L���V'��/�|h�_���gG,��G��:��!��6bq�M���ȉ�/�f�Q��3��`���yφ��oU>��5K��jJqF��|�!E��z^�A`u���D��K�v�	���М�v������\���U�g��Dcn�����͇���O�r���m������*t��O\I�uP����>�c�2�f��H�L 8L�O_��z�LD��Y_f�-�~�<��z�lW�_ �ΰ���-�m��c��޼�H�� ��F�p�����!�_N'�|����)۱�]�{���@gߴ�� L��eZVh_�E�f�v�R�ך��54����.o�2��nlC�!x�<3ſ�����_�u�@�=��<d,Q��̕5{�-݂��b��~$ǊGku���=��a��k���K���hD���~u�~�X6��/,���W�����k2��*�󟟃O#^B��\��K+��2���:��H���ilZ�;Ϟ�P-�ل�Z!F������6��S)l�kh"�@���J��B�� ����ԉOʠ��\�:cBXm��9��+��j=�uI2��W�i�C�g,�ɖ'B}o�)y��N,.; �5�*H���w�9�?�jyc�� W�����j����xB�0c�n�fJ70-�0C�`;�tNr 	�9��Us�_	WQ���zI�z�;�Ȁ(aL�7�՛6"���_��jR�'|�V���P"=�ĝ���ݯn�n�٣c���@%�k'Ywi��xa�NUYd��� �af��.G��g�|����R�`#)�xQB��OH�� e�(P���<�?��)T����� |�9�P1��ir�	��xhu�#t�10����@�����#�%���Z	i�3�B}�a�0�G���F��Ds�L�4�W�q��ig눈��&3�$�Χ�nZ�W���z�^W���8!8��\�t�/��߆Pβ�?h�1S�k�s���^ɾ�%��|�uZ"��C���N�q��P]��~�=�D�����|�/p�G�}����z��T��{��/J(
���H�s�)���24j��`���yI�щ�b�5 TԽ�����U���;������ב�i��>���4�w��R�������/q	��kC�^�N11��o�B�)K�|������q"��4؉Q7MK% %՗qU ��MҀv��3=��j&q�{���L�E����_��������WF���>HBW���T�'�x�Kg��I����P�S7*fg��*x�Z����svD5����nkw&���?�:��R~l}����^�����n2�����W&eޔ�xwuk]m�|�E'�6�:��EW<�$����8fW��
�j��A7ɤ�W2U��l���G�p�Q��	��
'[�Js��^1�`*�|>���|������5Czg�yo�cИ��x�T��m}���r�F�Q�V� �� s0�d;�癶V:ٻE0O��(�?'�2V5����ҵ��Q�R����;�EB?mV�X�6F t��J�y��1�e8uv�C덆��촶�Ç���\w���LQ��"��5p!v�u%�_r�UJU�/��=�+�������9(������F`�:"(��-2��T��P|r[U:&���1��T�;"�/�@W�O�bĎ_s~ll$�r'� 6�^��To�.�"�1��<'��nRFS3��lAp��wD��c6�*%�>�є�,O�a�ς���ʋwl�N9<�(�Ȼ�	�/���O��O+����)&i�hmb�KGG�>v�ن��V_�ϝKa/N6r-p�JBLz?<1�W�z1��{%���z ���dvh�x�5�Ǘ��a��2�[�w�J��4�+���H�n=�{g�+�����H��k��wH�1�BySw�PEo�@BH�9v_�'5��#B��<{�2O���[�����ʎ��QN+C!��"���݃��g�Η�Z�ޯ[W�kZcy��|;�1;	�;� T�忶�!���7��l�;%�rz����L�o�e$��sX7��s�zp�޴Q#J}��N%	pȵ�) �u3s�v�S����>�8i�].mdj�����RN�Q��������ֶ@ӭڬ_�T��[į��	��R9�˶�x����Е�1��H�#"���N���K+ؼR�R�����\no��x�o�i`�%Q��0�a$�x�H�H ��0n� �]�ѹ��7���5ɉ�R3�_��)�^�0��PXvj��
6����"��_zx���F/@�]*���/����n�EB=��V@bIO�!����԰��.�%��]�H#���;�S�����ֺg��OOO���f����	z/���S�&�/��)��h`9��1�w�k[���L�Qn˙�O�p���^�W���?�
�B�a\]�Zo ��ߪ%��j�
�c���L*э�k�?�v�MK&�,����f�xQ.�(%x��GP�q�T��n��H���L^&j�����k�+�L����Q�3W͟������n���H�ɕNw���(>{���"j��;��<Z�Q�ӑ~qb�%7%��P���@0�s���8��s0wF�h��F�E��i��}��uJ6^s�U�6���#n}�~���dÐ�X*�t7j���f��p����+�YpXC���I���E�p^`��IM���P�1nǛ��!���(��������m5�S~���Sr��6r!��H������D�tv�R:��tE��cl��T.��l�pz�<iI8G�j�Ș7f�d��L=���� L������ӡZ��\�$�[���9�X-Z���m�#2���8;���*Yjɥ&x%5�%U�K�u��J��^n_��Xp�W:�dg�]��*�j�'�[�G11���=i�x�f>���!da���%�*Y�Jn�wW�6DuH�_ׇ��������P�����H��?�w\>�N�7�@Mo�+��m��T1+*��SM�WĪ��`3
���	+/Q����!i�ۗ��xftH��SYՎ��g��9.<��M���.�WS>ҚYj�����K�Q�(�!?P%��<Q˷Y
m�}�^����\�z���Y�h�˖;��
I��ӿ��DGv��抦�	�%4�k��\l"8���x������S{�~y�W�p�Ȱ�;�Һ`.A�Sֈ���Q���~VC�A�R�0��Me*+�A8�̽ؓ�	��������{����4�=�i�).�4w� ���O���l�5�(�
Tye����qa��L�-�仨亻�a����=��i���#!�x�Q����j��y�z_7��ωȁ-Q��h�jU�vy�=��Y�"�O�)ۆ�E2������ßI��4��d�~}0V5��Á���|Ŕs+� Cn���O^8U����p�oL6
r��\	���C��Lͤ��lfT��Hߤ�{ v3
�*��?��o�e/ZMd"6o%W���W����VuK;�Ď�kr��J��;I��2~�ظ���B�fPui��)<9~ެc���$>J��0�MK^���s�8f�	ڰ����2�'jN�G��p�iT%���y�(��K^yr��C�F�X�M4���3��׏.�ey�4�q��zW�N�����D�?x�� ]��j�������!�.�=Oi�/
���(X7r�2zTV��h�=��VHMr���bx���nC����SmR#N����I!��bv�����RĨ����I�s��t�
4��2U2�ڄH�P�r��T> P6&�����q$���~�\WHE- �xe��)�����)P�,�F����RRhIf��&���X���u�H����#�tc���w��d�-x�.���5����gP��fP�"�A�.W���P0��׫�9h�[6�t�N��|�޾���U#lź��&O�$�i�l£�M럀>�N Q;`"xCѦC����(�k�TZ9�`��є(̢��8�i��a-)N�5�ub�#���݌u9�dY{b��@`lv,ocw%�$f�?8DU����,jǬ�U����#�׬X42�Pw*f�`�zy�n�ƺ�q4�������>��C��	���k�k�ͫ��R��� �1�BMd8�ig]5�-��܅����jޒ<.��T�{J����!4n��6�g\8����nڈ�溇S�	Pw�=WF9.�m��d�w�p�pmI�����ի\��i^��v��Ḱjy@�}�ҋ�&[U����<��'�-q�_�X���Į���o�
מo)���rb�[���a�l�'c�=㶭�������;�QO��&�H�����Ss�I�ՒU*�&99�����%1[�i��w0b4i2Y�|N195"C��c��kά����4��c��9����vp�.fv�*M����2��yD3�fhS�Zٷ������F��N��_P�I���?b�
�[����^"�os!�s� ˉR���2�̑u@�?`AJ�����XOn�yc�%�?��i� ��@�c�=MP���l:c\��@��N4 z� �h,7� r�;튤��^��h�ݨȡ�3[��Y׃6�"1{
��܉g�s��Q�4þnPҌ;9N��,mo� �V��ڞ��F�	=A�1P���6�9=W���m��wJ�@��W5;�jx�|]l՘��p��-��W6� 21D��NC�4?=�s�'~j�	�Hy�O#G'*��Ka�uX{�6���IkOJ��VD���v�m����\o���n��s��`����wՕ�k��!�uzr!�d�Oz� ����eVl�Ĭu;ξ/����f�hHY�am�c�b�T�r� ����oV[�mŁ��4:����h/W�#����6�o-*L��M~�*��{z�}_�E,�C�	���q�P�P�i��L�SPď'0.K�[8�*�[�;��1�~�O� �a�M��,f�	�>>LE�%o�Cc 1����ɚ�U����ߎ2� �89���Mid�餭L�BQr�����Q�3pSnQ����kNђ�x#`���k�ـev��?2~���$۴������!�gs��%�sɫo[g��=3��Г���]����u�YݱȟT�\D0B��K���q:r<�<�2U�,��;DlC<Ԑk�02�
_uޖF� ?����`�^䫷����ּ���/�c�s�`L2s����������-/��ԛۍ'I�:�8c%N�H�&ˠX�"눴�V�#�@H__Y�?$�A�}P��0�h&qfr��U���/9�bd�!���f��!�V���8��=� �,���k���/s��L�f?>=�6g�ֳ���`ŗ=6���|&��΋�	���[z���[m{2�*���ߟ��^,�u�}�@p�-���s���K�N����r#�i���a�A�U��|z��nU�"�2Oc��������ëQy%f+�¹e����? I�#�f����_1�j������;���MO�S�<��M���j����7�{s�����cN���z=�F~�և�-�����L\�����K不���4�.�a��:�$� 11�^���j�}��&�/h���N����I_J�=l����n(� �x��Zk����XPV�SΠ�f�-��<a�`�0�>��,(��Ƨ�X��X�0�JA�o�'���PC�fn��ք/�L�����߇UI�+�kKD"�P�)������5�5��'P5�#7�`s_�P���E��J�KF�2�����)�xPAFs�W�FҘ(�T_0�5���)Ad���(kX�@2=�-G%ͮ?��A[�Ҭ���P�"Q�C�P�E$���:6�c�S�"+T�6뾝�߃�Y�l'����	R��~��!<�l2@��>*�7����@��pr�2�;��B� �ZoS#��	;+���S�
�/���T���8����-�j�����L����ZRE؟���H<\��2��[������6|�P�+\:9�(q��(�i?������^�׾=G��b����|���2��m2��!��N'1[����Xt��	�$�5\b�<�ҰY�l�.rv1e������h��<�	��c��m��nk�֥i3��2��{�dVhV����{�*6S7m�������C�t�
$������~��=���} ��]�6H�c��3Pr-ڒA����J�g�j���ń�7`����7���v0�"�1a���fN=zl�)hK�+�@���M����>�.F>�K���J����'���I��՗��@�	�I�#D2��!ܮ�$��ja��r�ؚ���Ɥ��.'���#O��{*ǿh��?�e[�uБ�MGa=n��^gK>;/'w���ҳ�2Xv'5��ҕG7������k&J9�%��"։Ư�n��=/�|P	u�y�=!��.·��+%�W��U�����i��z�0kW�7�C�w�6���P�|!1ڞ� A����G��M~,F(p\�/ϓ�C�*���]�kʦN�BnѢ0Y��A��gx�%k~�a.��$��:+�e
Oz���of���j�Xپ��[�\����s��^�5]�n+�n���"a7vo�?9�I-��l�ȣ����4��t	����c����f]'�^l���ՙ�>���C�Ni�X�P1{�PO�^�d�"u������~�<!i���p�)�p@������-�2}����AƯ7��2��_!9��XO�@��D���i�������@�:ԩĊ��ӂ1�1���^���s��ޔ���<Q4��6�u4�v&�%��� �쁲:�")�I��k\>݈������%�;�Y�������-)+�:P��(E��/�͖�Z�yR���ww�E:{�,�#��e�Q��>��}뿟�� k���4�ͪS�ݹ&aKϳ$^�D:QHng���U���gߪ�0��Im��ݹ���\=S��f�a ��$�n*�Ⰼ�Q���"��2������k��&Goz��Ҧ�;4�6��b���ۻNf��P���/}v*�T����i �Vs�b��U 3���D�Z%Lqq;?������nE(�i��S�n��C�����%�	G%@����,�l�E`��c��}�Tץ)r��>`�+a�e3���*Й�?������g���b��(\N�6�5;5�n�Y�3��xC>{}K־¼;�<3����vF��7���NFC��C$} ��[&��".D��Q��֡Ph����-;.�9�Jf�U"vتS��w�p�c��Gr�ӱ�c�Þ����(���ܢ��kC�6�ю�ꮸ�����=,��H��H|��\�T̟lR��5��b=#,�Xx�a ˦�VJ�U�+jUm������3uE�Ik��������lB������s��U�[8VIr�W����@�Ft�'���, �@�:�Q)�u�߬�=�B���ؒ�H��@�;�NOM���e��=��~�u�D55���K@��~��w��h(֛ٟ�,ۈ�o���9,�Rٯ.��}
�LHd��x��I�^)t$(^�Ⱥ�y�����F��W��ۭ��t7�k�\H1���n��IS�k�xnS�	QU9�0�k��Ԅ9yF=��7�,��f�J�{��~|Ɇ:�F���z%"U�y���jj��Og���ʓw�$)6�fY |ukPD>�+u�'�BS�:�6x�!�=��,�w��6�nOV�!�Nm�=Rj.	�p�k���V	5��F:}ydz�a���c�+(�mm�NB��/ݸ���j���v<�)R���z�H�j�5�1{t��h`��=�[�X2��W3�^��ˋ�.���l��g�Xql0�Cę^������V�9�U͓�`'>��I����Ƚ_�F�Y׶��WQ��U��8��NE͂����&_��b�A��Ո��;�M�$&��9��\l�j�[���[�v;�X��8`�Rg��0�i��-��Bx����@�U�m�U����"SPQ��TXs{N���^�V����n hoL8n�����P��7�pR:�g�����򇶦a�M&���j�C��~f�V����yd�ԟ�B�3��������d<py�W�ڟ���Z)����g���h��ӄSqDy��d,^��a@Q+�]G�D���)V����<}���]G��OZ�BM���F�HDޘ�G�� WW��&�F���<�|W��&�?��~;KHCE������U���*��f�1q5x�h֯�U6[d���F�A��C�]�^aV���s~D#�J����ŉF奡�.��c"ط���*N�q^G��)NIű\�+�S�����@�Bz3��c�J^l�a��-�-����\|�\4�x�t˦C����5 ͱ��X���e�9^�IL��Q`�d(�Db��'=y($M�k�������e�Dl�v7=(�Z*jr��_�(u_������ɦ��S���oA0�)q�Vc��m�����u�.�����ܓg�ι����9�������O��K���J>SZ�10:��G]R�0q�+6���$:b3�n�I� o;�������G�d��Ȝ�R��\O�^���׮M��Yؚ�ϛx�`Lx�]0�ktqH��=RZ��c�צ��mc.hNs��*�!,c��{u��j�P���>M�J�����c�5Esv���[�@�È0�K�濓s��V ����@8Y�y$]�� 1��k+ڹ��Z;6<r|!KV܂m%m{Ch#69��`�&^�K�-��+�U
s��
��[}l$�����A�U{�J���Z�M�pSL�ЖQ_<�ҫ)�~sP�\�%�jϚ܀D:���Ff��Sz���,��`My7�B��P�/�:�B���m��p*�N���v��N�#1�ϴ6Ա��5�j)��~>�D<�$��	���A��'��D��^���ٷ�U項B ������ϰ�!��|$�15�O/lD+)�SV��f�����olV;:A�}�B�����
�O�������Є��ڢ���G�^�{�6~�IR����X���>{<5!F�2[I3^�'-��;G<��g	J]^1H��1���bv��VT?:<	��)Y�g��V�Y7��#���k���e��y��H6��c�=�]L���j���k������\�����(�	�Z�{�b�M˰9�K��ܔ�0�O�N�����*��t%��1���\$K�T ��
��l��j�eI����j��)7q1�2���eW7:�	/;�ősP�����D�G�¢c��|ד��Z�]�8�VŚ�o_��m*�T�|��$����U�38Fm���_Bv�A���r�qi�UH����0v2����V �)b6��\�f�G�!i�w�O�;����^����X0�{Hk�^,7��
�F���:3 �#��y�+=�iv�13�WU_"������z��Rd�T�q.=� �ߒ3�?�����'�3�Ez>�~8&��:[��>8��կPV��k���!�'c�M0��U�X)��p��#���=4�+�l:>��͍ B�ӆV�j�B�ϳ�g\�p �2p�J~T��L�T�w{gｩ0O�f@�C�$ޛ�g��݆1������d)�a��a��яsp�"�MX6�ф|�(�o�I��n&h�G10n�˫� ̬%�Rᶧ�����Л�����W}��IHr:�Gk�͗-���f <	f"֍+�o��S�f�ȑg{�M���p� �/[��C|��a��vH�X�t�9G@D�E��ټ830�q
�d�;\��q,L��N�B;��	=Y��@27L�|2��2�#���E�1���";��J�Zs�L��jg3�>G��cU�
$|�B��*;�ḣl<��&�i}s��݌)kP)�<#��ڮ�[��W���rpk(�$��7{/!��xq���@-y�zP[tty�S���ѰT	fÿ�<�DlW��4�{�;��$�H>��X�����þk4[9�yl��
����'�*��ywQ���I��/�����D����|�媃��'��D3:1�'�s�0´���6B8n�a[�X��wR�Dt�X�1�`w2c$f�����z&�{���-��y�-9{,�����Bڂțq��5h���\�\:����J�jlO��a�><�7�WݷM���%�=3����A=]�?�&0۝Zc*[L�U�����<�+��i���h�0LzU9.J��-59ʌ�݄��������\�WA��/��K0��RE��[M���X2��}goVьN�丗}l��g����" j�T�69��v6��kY�eM��%*��bmH3�ZT->�\q�rB�%7��=��Io"��X��U�AX�>������]F��?�v�τ�h�DN�?8U�q��mU��@II�guJm�}�Q�B��ؖ�k\P���:��������x5|����E�n��7iM.��T�4��y����H���Č/��Q���R� (�����<'��}�yTÛ��!+�������0��W"EÔ������n�	i �E������ճ��$�2�uF;ݵ����c�?����DbeG��އ$��Dz�B.���:��֡��6�
!ZNv?T&=@���bDJ��mI�V�]O��i�S��(��G�����k�v�S�"^��G������?,x���$���hs��v<	�	�
EuG��"���_l�^�e5z��~��0Lఴ�Q��Z3�L��U�o�j�9aD�
\{�ÄܿI)����!:�g:|�gx����,�o��v_<��D���c�P.�	�`08�FT���= �m�: �c+|��1�D!��/CTm_�H�F8��e�Z�,����?�Vv������凮\�-�oΑ��:2���Y�}_�+ E�+ܶ/�Z��Ney��У�(�=.6Y�	�����P�:��&����PL}v�6a�gT�pX|����jW̳��	��x}���~�!՜^|���[�<�Jo����bٯ�imOq��9x3vG:�S�E���g�ŕ�% �,�2B��H�6f�/��������G<ά���*��4�T�^��:�����*�⤷��Ӛ��i=���uAɝ�0ȉ����us��͗����C}�H�'ʄx�Q���}4��U�����ri���T-X��ۃ{�Ұ'�4�.�U�+��ti9��z�a/�UqLE��F�I$GƘH�wU`�.�7*n���ȡ��mdq��R�b��ob/y����/���v03��<���j6*��0���n�a�f%*��b�WvՌ��3��^z�ۆ�ɋ�ȧz�xR��m#o$�C@��"��\lz�4�]l'܎�y����������1mC=8�]�l�������g���љ����,U�K�u�� ���I	B)� ��\�'n�y�SՓ�M����r�q�9�dܺ��/`+j
�l_I����7�Y[���7t�
T
a32��%�dĴ��rɵ%Sp	X0�:�̌1���D����*k�K��t�%�T(ٛhW�#�lM�7�UZ@|�x���H�y[ ?�l�p�'q���W�]`��S�,�4����AZwx|fI��Npjp�HHEQ��FvT�mT���$��i�^}�!�ʳ?U�?�o+?�ɅKGH�ng���U���ꁁ��~ʟ��,E�`�h�u��D՛r!�bGq�K��1y�5�Tv$�yI{.h!UR+)����$����S_�~��=��)���� �f[��J�k���}'�k�eS���9n��*���5~�^�GA��H& i^�6���T8x��'�(\�ZqW��|f ��-����8:˟(����X���Cr�j���*ىf��R��M�k�,�sl,������+��¨^&a�D&��B��`A@�����yI>,��{�Jسj�#�7�E�;���k�<�f����xzh�U�G�I#���e/�yة��Sk�+Кl	r��Z�n��laf��1n`;��p�����?�ٸ&1j
�;T���bpu8�d[�t�+�gL7��q�y���S�T+��y������δ�ٴl��Z�p��B��yZoV�<n\�Nî�^��0n,�[�������S.~KuAh�y5Hd*��_���@�Au~넍��I�悱��ФF3޶lѩy> v�.�"#�����ѧΙr!�5@/�
楗��m��s<��r��2�\�?<r�����Ý��̸?z9���g�C�z���e�B��샳�\��o��3�]jZ�)@O�V��x�j&8��`��͊7�?OG��'��a����m��$�o��guV�%���
o�AIs��aWV"`�K�]n�5)+NY)���μWSK�Ρ���E�{��e��-I�2y�h�{^!�,�"η��i�\熡[#S�5M=�L�&0A����,;�Z�TT��ڏu��j��H�x��ӈ�LdV+�bo�]pso�t)Df�5���M�w���FZ�$���/�ȉ$�TJ��q�2����~����5I&��vN���_HU6`�|�{��t�8��J�Zơ��qQ�#e�ؔG�����.OE�ش�/�&�5�\8@����N�-D�y �odt�ی�$:E�o���G(�+-õ�q\\ Ǡ� ���~�X\FW�²9�͠�+��bM1f���vZ�<�"��fr�����*c@Xb��#�ix����ފ����n�}*ծ��+�9�	��3��d�)�VQR. S��EP1�д^4�:�R&�����HF2ţ+$����W{����Â��*� ��-�[ϓ�'V��u��aD�d���b�7ۢ����u�����2�
>�2ZY���f��9�Ћ�-iS�	������q�v��Fr5�Z�� ���$�?�0�)p����F����$J�O�l� ���g6���D�'�L�Á(b&'���j����T�c#����s�A�G?.���9��O��_+V�4��T��*+�q�F2���+�4W?{����;�9�$-H�U@?�]�'�DY��4w뫉��q��9���4�ql��uMoP�}Ӿo�8E�9�cr�Q5݈��s��Y�O͝%�n�K�^ y�������>��Q��L��n�Uf���t�2�%�<ڨ��Fܒu�~4ˁ��s:��ouO�?�>)6��݀��������(���U3���]`P���B��s��U6��6q%���'���E���"���ߜ'8+M?jT��î�7��Ej؛�
ՙNqi*�F�0�3�ډ���F�TI*˺Z��0ŗdUSM0�gm���0�Y)�=D0�c����
m���U�9�pfH�6R_�r �e?7�����S<���ځ�m�\�
��x��|������1�Q��J�a�����י��?�|o�\ď�M�]���[��"ڥ	���]-s
[ȰT�4������ku��yӑ�yM!��[�1�Cx�^*�Ua+߆��ġ��E�����P1@#	�N�Ͻ|"���_�3�t�"^�*j�_�⒥��*2Z?��� �y�şp�%>ȯ����/��̨޾���N*��[��gɼX�s5�(Y�=n�B�?Z�ֻ�����q��ض���k�;s�9T��N�
6�}钐�%m�N
+��r*a��B���f�֖ԏ=WP]��K�Y�:�0hz��$ g��ظ�SU���� �;(d�=������h�޶�s�~TCy	4c[�q��n�(������p�КG�U��,c�K:lq�_��l����UX@�1�f+,D_�x���I��F�fo7"a8����Rrs`���sŧ���
��D�b���C��:T!f5a_������JhZ�ȉp�͍1v�5�;R/U�Wu��&��:/��{���9 Yn}�w���yЭ�*��UoM z�z����������z��_�'n�������[��=��ecI��|"�m{ۊ���wL=��OK�/n���=l����՘ǄP��3��s��Gt��@�L�3P!��`A�����V��.�ܫ���+��A_�k�� �p�*��*�rSI��i����,�ȼoS�VЪ1��t����\p2+R�V�RW�h�D�❵ط�F�)�'˫�)�µ7�$_�wL�R���0>V� ԇ���O�w3� ��F`b�ؖ���[��D=�j6{��B��]�%�I2e��ߡ��
�2B���v�r�j�VW�v/��bc������-0c� zT(a�4"~R�i�y�?�F�>}��_�2������ܡ���O:�Ñ��:���p�Ⱦ���hs+�B�S/F�6kIQ@RbB��n?-޶�*��T́�;��=�'sx0{���4��\*���B/�8԰���OY�'Al�¦�Q'��b����+�J���<�*i�j�,�D���&��6e�s� $�8��V6?��u�.�&��\�&D���#C��"���2�ܵ�L:�f V��G ����YT/~�>��Y��G����Q&�t�^N�%f%� h�����ɲ����%4�LIe�#��)���˾CP��`�͕������$m�U��>Gwv:�H֗9�1�%�m�\�.���r�r����k���o6*�jsFucq�kd�)a.=xm��:�m~��וr�� ���kM��r��x1ą%B?��Oj}���9S
��
�I�m� |�g�'.yd��ێ}�!�v,`x�O��A�	I_m_B�E�x@;�g0L^M�B�-q��U��2s��]xb�ց|T>��jyf§�~�n/�����B��V��ǢӠ�ۘ���?�3�����[5����F��3�3�A�V�AV�F�M氕�a����	�'O�Ci��c}��P.��|�Va���e�Ӕ�<g��$ag�4)�!�,��g���ݝl?ZZ�Oe�"���@�0{19�/{�����2a������찾�m�f� ��h����ۻf�6EĽ�v����@l	JyI��J��>&�;ɛ��Y^� u5mQ7Z[�J�\�t�Ϝۀ���c̮j�3o�W�<�Lv;?w�X�C��U���V�ۂW-���͕����[�iNk�������9�<�
%d�5�`"7�j��yȋo��/���e�C�:̕��~�������N������د������p���F5�D\��=9M�z��Pzx}|G\tv�]|��6�>�- �$.�3nz'Ϧ������p	�;��,UK�n���Wp<�+���>��06�����L�hU�XO/��{�<�Gĩh�3ԥ�^��q�[��P+�����/R�h��O=8e�v�����q)n؋AVN��=
`O�O�?@�K��"Lo>e���rx"��ҙ�d��Ȕ����f�%��L�6lS���,�;R�\q��3�1V@�P#=�nn.CܢO����v��a��Ϙ�V�a�1�gjr�fi� Se��1�K�Δ���t�}0��1T>�m5^ �����=S����Gś,ũ�@d��~�W����r,Br�R�\���_Z w���;�V��ɭ���'��>V�I�EmTmy���
������8�G�ܜ|��ӱ<��.�G�N�`/q<���/~����4��� �إ��3꫕V�Q��i��
�4A����g����&�W��t��)��B,9�C+*�9ʺ ]���	E�����8:�x"%���E,p�f�*�Ug��Bw��сA��ʕ����8Ѯ�xgvm|imc}(���Yp�)��/vh�`.��]�n�+���%���'�b6����?{�h?��aq�
���3���ů*�n/0�>�V�2lvQj�ν<�k�ň��&[I����g�#:�a�G$��m�.`dİ ��(Z4
� m����׏��1_y���z�]��~Z�1�Xoc��$QY�J-m���WY��2rQ'�,�ho��������ӈ�_�c6i~=��E�����nX���r��d8���Q��!���QW1`Ag:�@f�jM;��_~^�b]�
G=���k�����X�<�@ʹ�i�p�k$%@��E���9˙RAm�Xo?��<���}5%��3�_6L����4�<V���=T�2zO;�+��_~��? ����5�]@E���(�﵁],w}�*�|�xY;�ޱ���\��X
m��j�����h����D���,��pA�R��T,�@�����}D��m7	�:��C1�
��HX� h�4G6�m�3��D�>b�8�R��")=�f�wျ�.(ȇ�~�IsP��4g�LJף��&ѕG��ˇ������=��w6���Z��ņ�A�W۴V,Љ$�Rw�o\v�ȥ�U�[ţ�"'�-�J��ho�8�ܬ|�'h�����`�B�f!=$�+G3��A,�4䏒R�n��v
�Tz��:Iҙc�1���?'y+6����n�>\�N����:<�����a�M�u8,�y&������譈��/c���:~4�&ɋ�21@b���/�o��J!`�Z4|Z��|���H��{��D��@{��%�x2�i�>��&��ܲ`	mM��7���1�]�8�p7���Z�-�1J*bK/�^�@<aPh7U RE@�O�gl��n?}ՙf��+�����g����ۙ�x�x�x�����n�ӎx�>\�z����_'?�7����������6����%0]�������%KkZn�uR�q(ݢ���<܍��!��}1�#4��g~�i~��'�ர��:��ﾴ��1���~���:��
�Z�q��&���g?>e!h��2��+�qaF��_�Kk%�$,1��0E�r�$1��5[��rV�re��S/9���� �eQ��U�#1��a�<|�=6���|]���d��?\EE��'N��Y�Eӛc��H�fL~:a�A�G+�y\�s���*F ٦�"T{��C�E���'[J���� ѱJo6��A됽v)�*$0� ��pq���.'��C�wf?A*�m�k��@��j[�X-���������r�Q���*��!~g��f1�P.1�<蟋��`�܉�.��ߗ�J|���6]"�*��r����(��6�g����I��z-�X��U<��?Ù��)Q��Z5=�/X;wL�����:��'��X�Y����"bݎ�%���1s͗��F��������[�����#
���R���⤀s̕"� �(�&p`����ޓ�v9]8x݋��������2�^Ho�D�����}��@�DMB%w�2@$�o7>S"� �]u2N����&pܑf�QϬ�(��'�y�6��#����
�:$0`��4)N9 I���-��K�Rٷe��	b��]���on5�Mn�e���x��.>�3Ҳ���p�_�Tsc����K�<���C(��O��t&�!�������.tEs|S��������
��R�p�$�w}�kiO�)|�9D�L�W����b�eGL�oަ��~�����l��F]'ݦ�q8����_<}����RM�g���ߖD��Z*M� �:�ٴ�<�������mۅm
*o4���Tt���PV��Eg촦y�<�g��};�e�D��WYB��#G�2a��Z$w�����Kr:,�x�����s�I���#�O���9Mv�Yۗ1�Ğ�y{ � y�KT�|��u��>F���F�,����pI\n�.��2:	�R��⡐��ӝ4���SI��ɦ+H.\�ڙ'j��^����y��7�G������E�|h�i 5'�mB��%,�L�����k��A-������G\�	��Fx��.iAR:��Q$�N,ψ}�?���=@=��2�C�XFM�������;�?���&��#��[%�#�b̾0�D,49��	v��k�u_[�M.��q\��fzê?=#.�;�1�s��7�<��ޮK(|v�A�jWh̀�p"Xd���϶���w�m�N�Ru<xŕ������	e����Y�B��4��%8�*J����FI���B$�B�	P��s{��h|)o�61����X��W�@�2lV�ʣ"��/�Q�t�W~��U������\�q����:���F�I�EjGt�VP��e>ʨ�Cj0h?����Ќ��!{��9�m<f;b�8#!皪��s ���#~�=^AU��Æ����y/ �,bŮ��l9�Ia��ǂ1�)ڀ`�j7���1u����$�Cj��$��S�Ɛ,CQW����-2�f:��1c��5���ST�'��+h��ޙ�)k�U���e�)�Uy��&��I"
nCF��UՃ`@�I숫1�2��Y ��C���"�h^�]Y[�?�Jǖ��0�=���C��Na��y�wo�0��h��Ub����@=:�WQ�E�0f�V�n�3��o�_9Ǘ��x���5w��8�	.���X�)�~&B��`��jy�Q�����,*���Bƺ��0r�Zz���|ɚܻ׭�D�����je���K�n�����9.ߧ{K� P*���X=�?��Z� ��V�w2n݀�54����(�aoTo�篎�[Jӌ6�@	���9�@��!Ž#/�	�I���NN�-:��M���� t �+�v�=�o�M����k��[`@�q��2*��x��tO)���؏.�����$���T��9͡y�f�Q� c.�&�����*Z�
��O��v��|� �̶�"d�w|,��u<xхvjVإS���S�S7콹�6�7�ͥ�<*:uI&{A��S������%=�6@�R1���m$���j�0��U�"���L� ��o�
�4&������Ƣ�=tX�z�=?��a�Gl�j�]{��ns�񐊝I�md��m�}�+ʴG���yX��Ly1�B]�r>�ȹP��c��>�L�<�Z����GZc���G��h�-G��/��c��x[q(Y��mh>$7-�|H��	��. �}sF���h�r/|\J�|_�����@�\7H�g�||%���\(ݶ ?RL�F�'nܻ����u�qj�XM:����٩��*��!y�H��&�Z���i��^�㸙�y;��B���ECÄ�8�2.j�J����d/��0u.�	�;����ƣ���(M0,���0Yv����(�n!�񟠁z��^uX,�R�x�a?������
�;rS}\<k��j���K�kg�Y�����nmn.��9ƈ�K���-~<����-,+��qJ��S$�G.���7��)V�~�h=س����_4���'�g;�f����#�p�U�g��Y�yh .���BiI6�a�����¬8S��/��r4N�*_C��Nq�����V�G=}f�G7����%�G��<��|�g+	f�*l-8WV#cz�5/0յO??;i�u����@I��ONl�"u�����l?����{�j��/���a�׊`��qޞ�c��5������*&C���;��e�],"B!T�ɝ�t���\��486���c��G�`}M�N�^�	��y9\(�pm���s���������3��ū��\V���A���:��V>�S�ñz��,��j%����X'�0mp,�~�A�KP�WlMAW���2�E0�c�s]�DAw�M4���Kt��4A��M 1Fl��q��a�_��`�s�(N���	ކ����w5�?�}y��B2�Ɵ~G�Mi"(ua7&_?�l�X�;i�~��׿����bJ�����7)3���2\�<8�����0��5P� &���k0��������h����·�<sG;���j�C�c��ďHs�Et�,۹G,��~��`�4��y�\v���_ aݼF�ҳ6O>��]�r�%;�Jv�!Z�"�,�f����,G�rX �[}��氇�C�@ &UzPsP�ȹ��vlhǳ%O� h��y�4(g2_�_oO�Ke��P�(*�2W�K����H��:�-�����X����w��T��օ�(G?Lr]un	�1f�VLE��p��{]ӿ�$�y�t!����U���A �B�u*�<�<�[�zL���ۥ.��:�]�{%ZL ��rsG�F�)����W�`�g��qj�)���%��d�4�����9_�-'q		҉���SJ%��;0<E^4��2n��C��v�.���u��l>�~(o ��;W�V�K/ڡ�ا�o�̱T�9���� ��}��`�2۩F�t[n��zM���V˙td�+��IK$�/p"T��:��j�N>�6� �z�v�`�t�X$��n��*�6�r~>v�KD�,^G�ӫ�|���\n�4�쾵U�W��9�!9�r���
oI�m-m�+H��D�W-������J|�z�����~�NS�TF4~�fs�b��9����Q
��]y`XA,g`-]`(4�����u��P)���=K��� .Q>'R}��w��ga�%�zi�A�.٪þ:�7֯�yl�ݥ�����-�U��x5�Y`{PO@�Е�ŵ� 0r��r��w^Gbdۦ�ye�Q��r~��u���ě����<�p,?RaM��l1�V��9�lCc�ʔ0�;/��,W�v�}��/9�$����8��* X��oԅԸq�*�{��-y|-����帚�2� h&f�ōH�e�Z>�\P#�ۦ��D;<}lfO�񸱆v�ؓY!@��|ի� Հ�ڒ���� ���e�_���t���oQ%����6�KoR�v�S�g��/�)<��W�y�H� ���c]�^a�T/�����c7�~�cHWrNڸf��!pc�uHd"�>�R	��py���������E����-�]�����Io���D#"�d�aCP������/׫�D��ȭ2͌�_xA^.��#�yo�Qm*�Ӗ��ٕ�rG����BI����$��O3���q=L��"oP�T`�F���m��a���m�����V�ڇ~:C��#�p�1G�h�I�-�:��9�K�H4��¯�E�@GI��Z����l"T���u��{�n�]ԣ�c���hr�r�"il<c���S0e�tg/GY�w>��/��ɗ��WO�G�v0�(�'vC2��[���g����
�*���(�m�&����Q�~-y����U��W�s~��@'��ʍ���՜x����|�[I���W��x�tƳ&~���Zh�����T0�ņ�����H��*,n���H(�xԦ���3��h@�����z�Қ���ڿ�<��Ӫ�4y(�W_RHZ�����e��$ˆqtq�M��;����zr���ѩ]�J`�	9�_e"�gSZOP2�)�b�uߕ�F
c�Ukb邛*W�3��;�E�vfOk�p�ù��);�h��fx���Q>�SX_�6Cޕ��>����hB6���;�L���
����~�7�B3���~q���S�)Dg�4�r�W]�����t��*�j��nߌ���AR�&��p��?�"��+[��f� �pe��3۱'�5s��ڂ���^�v�x�F4&t�ؗ7�A$Ӫ/f0��� ���SbBK�f~��;F?�#��D8�Β(��6��M�fe���ϡ�
��)�:6=����E�I��(0���ʁe$)�\��%|�w�z�o;�J����œ 9- �(�@X8�G�'�J�~��)2Lj��WoV��P{S��C m��m�b�T�^�}�t?u�J��I��3���뤭�?�V�����׈Iv���C�%�i����   ��V^M�I��U1=.��q*��B��C��A^-U�{������W�?w�q i"QPR��3{�$�]b	�O3B�C*u��ںP�%I׳_U���N�!v|�*���y���_I�S�����ɺEZn{/��0�K� +�I���E����L�"��K�+�2����ѐ�����)�
�LC�p�Rء�#�|i����L!��q&��EO��}8I�ܸg�kU��@>���jh��"�7�f,U��Z�RS`6':jѯ k�l]^���\�iΫ#��#$�f���/nv������� �:W�#���� �37���~���O:�# �s�<�*��p󾎪!6f�?�a��n��He�q1��^�Ii�dR��S�D���� �H��NkPxl���<�M��W.r�x#���t5������ Xf%���4[ܒ����A��X[ �Wxj�M�˟� �-p�;����)tA���@���):�Tq�c�T��/qD/��7z��Bk�R{s��M��]���oW��%Ķ̽���ɔ��#j��{P��"�"�ƅ��)�(rIx����쥷���m��O*��08�zQADLx��!'�iOi@ܝ�T���2�1��^�a]R3<Wf�a���e<���/�nu^6�25����p��c����vcF5���N1�J�H�V����Hx)4�4�k_M�a��l����h��P���l�tDg{0ti�5G��)k8���Q4���q��ENZ��`����Wj�Ap���� P�I��U�L�������0�x�e# h�vB}D&��L)\w�#;�:_�m^����̫��M#i53Yp��[���QI(k�$ZfuU��ꊜ��#�8�/����#m��꯼�u�ZA(����n�i�y�/�dx�ߵ4*��	nY�	Jǥ}	�,�u�8Ib����t�)Y��x�]!����KCo��j^҈��C x����wGi��J�"�B�N#���b�AB��8�]�=�G#�=SW�S���u���x���ڋp3��݈$�k�u�q;K�
!ߏ���� z���+�d�d5"���ik�.�0�0�b���Fo�:��D��%a��0ݮ�v���DB١����������Ni���\�̆�9����f�K�gF7d(��>c��p�#����k��_z��:���G�5��`i�����.�=�eJ������Lm�"�E��\�]�ߒ�V�0U��NC�x~8�4?�'2,�-��~�����>H��B(��gA�"]`�[]��V�4�A�M��4�G�m%S8�6�,�d�~-�I�Ӻ�"+j��Q�`e��`^fޯ��;��Ƣ�6/��>����$�nq`��8��yvb���F-pK
����ذ�6��A@�`[)��1��$����h�7g�3bO�~�'*G�z���R�'I���W�a�4�SS	���=����� jK����*@Q�����x���w�j�e�f�}�Om�b{�l:����dڟ�/�n�C��*k*RC��dΆV���~��������o��~]��3Q�bö�w�XQ�?s*�[<{T�B/K�#m�G�#V�Ӷ-�N=�.�i��G�����}� eI��G�����;��#���-/g�E��
	��/�v��hN��M@�L���%A�t�3��%� ��x��5`�i�Ik�����$�c.�����P�����M��Y�a�r~�"r�33~�jEڢ�Mvi�'E��=����U)~��p�	5i1��� �C�g4�'vKuDD��s�Q�X�N���� ��y@Ϡ�Jϐ':d�������!��1�����zB|̧�~"̑���n���c��C�s����5�%�ұ`�l����F�N������[��ָ:v�ݜކ�e`�}'!���$JG ��Y<�W*%� 8h�B�O��xT.lV̨��X� rZy���
�@	�B*,�q/�:����en�R3нl\kgBh#z��<H�0�����ʦ��=O��Y<j�5�a��ko���::�Ev`$�~�^T$ڋ ���V��pgp��'�iꆽ�#�fo�0c���DF3L����G��$��T���PJT�d?�`/Ű�o1�a	Ts�mQ���pх*5U)�ё�u����m1bB��U�U��p>C�DO��N��y�&e
�ń�åh�˝�΃��aj3U!�=�?��H���щ�Ļ�}�|�Uu���4S�)Ef�:����4���=c��n�o�M���S
��x�J�����iXxy���+O4PE�"õ�<VS���q��X9.�<u5~~\l���~�M��&S�W��fV��3i��I�2���5!�ό�')&����	JP�wB*iQM���/��:s�y�%f켒����EN�i3Y��`z�$�}�@m�<B�xȈ8&�IRP��M<zRЊ��S�C!��������C�)?%�h�A���;@QW���M�_�=��`��!ϟ�����}� �q���0!D�E6k�O�pW�������]6s���Y�2K�O�	�o�Bb��:Row
/�w�]?5e�o�9�-�! �`䁵b-p̭0\Ϯo�h��Ò�EP�7��5&�ǫ�@>>�t��f	���?U.��:�{�*ND!뗯q}�9w���÷�ɡMa�𚑂��XU�d�7I��_���C���"�~G	���;�BR$��S�f�B���+6g�a�� ��k0�jn}ȯ�ᚱX䀿f�MMRA��;�Un�ܹO��C)<KPߜ2�A��e*�T*�֮h�� M��],>% f���]��p>�i�츤�M�@������Zz��S	��3i)��$�-B�(����({�˚�8F.h?�A�DN�z�:ʬ ��b��L��*�|:�yS�ü[��KV�5�oq�e�l/��$���QV�Ƌ$�m|͛�z�#U
S�f�y���y;)��|���d�I�d�*0����b��}�c+��XIŴ�"Ԝ���-l���(f���5ѱ�䲶�RsS����W�( adHS۵�'9�4^[Y���a}=��
FD�В����%C��j��I(e.��U&B�C;�"�L�+8p�%�Ax���/*b�n�f9�pªq�
��^{�>�$xi�s�:���IŨWZ�ނ�L����yߜB7�i���8��^l9�� �'�5�_g4�q_�l�Q�����ԭ��D(~�TM�P�eǴGig�1��1�Cs|�v}�J�HM��P��>���^B���<����
:�|�Gu(P>�'�q$��nM�Z.W.�������{�(�!��	�<p1�_z�1�q���c{.J\�l,_�񟶘�S�s�&#�����k�w��T��L�q J�a\(X�m�^�o�kI�t�;qe�t�N�u\�a�ɹ�M��٢��G��o坁= �`p_,Y��l�x�����������mH��������S�,�~�+oD������d&F�&w��]՚B�䱆�q����I�J�A'�^��C���ZD�Gt�\(
Q�K�Ɵ�;�� Q+�5��+	b̧4?��%���l]�S��ς�j
R�83b����*߄����V���k��ɡ���ʻW��s���)�E�ryh4�߸�|\7���A���%K01 S�S,<[�_��v~��1/^\���b��z���p��q���k���F�p�����V������3��qϛ��-܎���4�
ж��oD�:��9^������7�M}��l���r���^d�q]�e?/ n���	 �����h�~�b�O��m�%NY
��c��Z_��@s3�y����� �zG��^<<���fv�ۍ�mA�X|�blb��w�N�5�����������7���о��TB���=v������rIޤ��Z�$�_!� ��6|@�I�k1E�]��ry�Q�G��i`A/�z}����}��8�P��v�(�o�*�^]�򂺢�Z�5:	SD��f�%��
�C�UxZ���	̖C�nN�����q�赸��{0�Ol�Z6���ŅɗC��tuE�\�����W(1gZ1�����.�A�4�v��i�">t�$�n�f�
w��7�;Pc�.��/�g�����"�-�{աbF@L�I��h�i��QJ�GU.n6W����p��n�խ�}4�Gye���a���H���;]x�ԗ��i�m۫M:p�p� ���������t�ϒ����?��q�ؽ6S��P'^N��XXC8��|���fz��B��o�G����J�)��K1
���f*2�P�������;
������#�*=���F`a�<��Կ��"2�?hI}'H^�=�paN�'yH'�Fʥ�B9an�d��S�Z�s�]��tCl�{�:���+V��"��m��u4���@��;�̿} [���z�9+'�T�S4U�lP#.O`���d4͵���"Rx"*ЍI�R�\G÷�4&e���?��GC�s�T� 2	�Z��
�*AV�:�k1��s_��{��g��bC���~U.7W6������r]�kI�qH��l&��[�DܻHz9�J�\{���VRg��H��L�ƃ/�R��L3�X���mX� �Ȉ��m44�C��|Pc�'���4@RTФR�����|���^�!�x4	(5f 0"���5-y���	��[�cK8Y���}GіB�&?*������L��āBií�����!�U`�(�:��z�Ǧsr���W� �xoj��17��֏�)c��Ulϙ�h�+�e����\�~7�ð*\�"d�	�Kh���[� .���\��J�;��*}��Z���ӬqY��or� �2��_m���$��]�P�_+A���E�8��j�_���F���Ψh&m�[�,Y��������W35WG[M�����k4@�N���ҷ��e�
.���խ��Y���{
�D���5ps3:dm�"L����_�A�p�kPF	�A������Պ �:cEpq9���"�u��`�voA��K#�x"��;�<9�É��1���(�?W�'g1��?N@`Y�p�`�_�PΤ	S���|��U�ZBS;]p��ͦ(�o(ŉ���5^�i�<U�}��;69��:;S�-j�"��O�ӄ$uK���V��@=����ӊ��b��u��J���B;��wG��u��z1d���֩�'k�y9�/-�R�v}��[�N㟹�:��~ob	�S�P��T�] �k몲�q���h�8XR�\���'����őe����{�ǰfބ$A��y�~3G�>Q�
6��xڶ�HZ74������3��+&�!
�'�L����D.�������?,���w�/�U������p��_x-�ǡ�d92���48���E��Lu�V
�_�*��%�]�O��-���P�%�G>�*
����ϡ��~�3�N����>d�0j�w�-��+~��1��<�x���Ĝ��ɍdm/�5},T"���Tat�;�>��+��-��Hf��߾a}3!�Ĝ�S�v��O�^� ��-��F��4���4c�0t������K(�J������g��@_:/�m�N"�;CȽ��PxKy��ϥ�v?�6����u��1j����z�hB��l�|p�v�k�vMiD"gJw�s�$-����r��`�Q�(&�ڶW��)a�������D�q�X=�,���?l��ӑ?j4z	�Cj�=��p��/����Er"�۱:�>��r��ڕ�x@��lp��\�r���i���p�$��n���ȽR�HC�Es�q�B���(��>�����M+r�lј=U�W��6�����1��1*`�5��g�T1D&�>�^�I"UX�-*�G�>�,ܗ�}�����8$�(F�u��L����]�.
�v[�/�B�^pX��R�뛘�hAm�:��=�7��������fMM�����1�8C�l&�I��x���*	�F~�;�	q¼��5��Ӹ�d@v�q���	 ƛ�-
T�V�A�e�F�ǡ�K��I}�Hܺ冁pԔC�K=��"�ߍ�LO&�}*� �8Ưp��M���\�'��b�(L2C$UW�;�/���U�݄��Q́���#q���6�/q2� �E��Tce
s�������\��&&a<��8��
� EC�$b��)�����;���頢�?BR��ԘL[��g���$s�&'�ZVre��?�z�i����
Y���2�!:�F��޳OLJ�!sL&�n>!|gw���(�����v��]>œ��M��cO��95���<�3�����8�S�_����+�������;�I:P���39yD�x�o%�		�=���6�H�Ah{��8jwGs���d<Ҏ|t7��E=��Y�N���w�|h�C����G�v������/��!�c��� eK�<+��0�]s{w΅],�h�L�Y �"����hc�j��1�H�~�E��vĔ>�>��ۻ.?����L�E�.�t�[���p��m����nd?<��!��jq ���E� ���x�<�$��׳m��h��Tr�D��]�"�A��#�ٶ�Aܮ�	��,뫁��}�\�
)Y�N=�QH��iEBBJ�5��e��SNmw�D
/W��%��j��ܱ�p�W]Co�w���ʏ�_�u*�?g;��z�=�&�����ܣ5Z�Qwdy��S�<�*Z�c��KLՊ_�w��k�����?�f#��Z����~�x�1x"��eO0�c��Q7��e�Y���ek-wf�YȃY> �V�J��^5���؃�,�lr�uڛ����@1/R��\.ԫ���\�Y�|��/�ϡК7�Iȸ���g4D����ݢME����I�?9�X��4�~���
�D̢#��(?[\UAτi��"��N�J�؁,i}�+*Ga�ƫ����j����À|붪	��S��JU1݅0Z�o`QU�`T�e����:D�d>3�|nBRl�� �W�q�p\i����j"��C�W�(K�	��h��*��*�GZ�kb�!�a�+���	S���]� �u��P������!�9H�������V�75t�@�(	AP}.a����"1��wK���YH]W(m�d����S��xߩ�y�Fnn�m�n��Y6��}��/wgK�@�v¡h��A�XmKM�6��}�u=�$�2F'��^�=_�e�H����	l��֪����X�>W.���8{e���AQ�c�?>k���؃BB��t5��a�.a��Z��t�Pd�Q	Vs�Z'>��BZ��o�Ӽ,3�_��/f�'�k���?"(��6��c�U�1c�K�+���L-�Z���*<��r�MV@�o˺J�bQ:�u�W%�@>g���K��w[�EZ-&���,��/�<�v�6����_Wo�{������c�Sk |,�D\�4V���m5��HmA/�R��1�$7.=>H�w��[�\�M�)���9�Q3�BY��Ŀ�v�]�������C����2���7�����08��U_��5�v�����OI%-o0`!�w(e[�>�s�8�l���6���J��I�Y��V�+�����u{Z��tS�K�E��Q=2�����ˎ��r��xrNC]~���Cޙ���䗄0H��;/.M�]bMo^�� ����>��-�M�5�'��6�@�Qp�ͷw٥�� :?���/�ǀ�0��8W�I.���'�"e�wӴ코?�����*���C%P"���s���O����(��y�[�a��$K,K�p�n�f�O|�0d�/-0�fqŧ=��T��{�^�h�w+�3jmQ���8���|ы��v�k�"G��@��-�&+0'f�,4*��œ�?^�N/Râ{��h�s�Y4z:�Ce���nש�,k�]��ދX��봸�e�������L������Zje(%�ߨ�PV��뙩�4i�t�����  M��!p�{k��3�H�n��<r�/d��bOd��ԁu�+�=$F�)��4��o��Ǫ��^�\�C=B� �-�<��̾����>�կl7N�(�Ⱦ�wN����
�Q�E��ҋ&��n� �r�Z�B��F����?Qy���wW+��9I��|�cp6�h����3�����:@�;�H'g".q�Y��f�ڊ�����l�^���z�6�ŝ2�&rA�e��
�i�*��� �^n<γ�4`��J��)�[ ��DML��U� ����שZsg��)���zW��7���̒,�̩t5�"M���Us
�W+��4���r�HY�VO)xh��ۉ�V�-�N�M��������J������:�j�#�dl2�9a[�:� �"qN����V��Cx�N	px��Z�vD�NDSs$�</
C��:���!��|�Y��wfV*����uҋ����-�	A*S�V_P릇�J��Z��{���@���(���1��7GU�&U�v����W����4;�+- ���u;t�[�R�қq�l��=�jT�em+�og�G��̎�g6Ԫ��-oOƭ�A��?�n�F��H'�m:Lj�x�0��XI'�� �ս�y̆��󨲵��OQ�R%ɲ�෻ψ����:�Op�Y�r�Y���G�(���y��(aBC�.���Q�R���!NZh�.�U9�&-)�tyg�����b�Dp���v��$qH�j�v�4oX@�Ku��v�4�夼�K_L.����B>�� ��/��2�R��G&��n��)�)>�.^�w����i�op~�K�(6x�ͮ��v�Mve��1�=|�Hu��(g��\���7��ہ�����lY����{����K,�m3���q��A�o��BZ�ѐE���N�"�?��dՊ�����F���/\�S��M�$���Ա#�{��)�.Vh��*����7�)��/p����iQLǙ�F��4<J���)nP�:i_ ��C�MR���9oXa�Ѽ������Q��:(=�]��2�[����M	[a샀^�����ps��6��d��QV_�[��VR�g~�ه��S�Ї�����`��z�g7��I]�������2�MJ�?Ō���x˨��{�u6�
}B����t=x ���`����X�J��i)@ۂM飑#~���vipi�lX=~X�Y֐`dBbH'��F��g9k��7`�Վy>��T`Ʃ�ć�-z�%(�s�U6ҿMC@���a��� C�El�ʋKrRI3O�L�a��ه�<IK��ֵ`+�C�0�]�з��/�����1�˯R�"�m��8��X,�V�ĆF��o���Oa����r�N��W�b���e����ǔ�����c��v/Aţ.����=��������fbIOo!g�c߲�1����I����{rLVA^��C�P���Vq�K��Jb��-�wmCl�#a�n�&7��RP=]��+VJN�c�x4��s��sm�+xH�c�&]ܺ��m�g�[�����g�G3�Y{=�fY��rr�|��(����{��`	d��j&��Kg�
�2̓t�jw�o^�5�v�Mΐw~�
��Z��0F88�!� b�qd�*��N+"�h��s����Q�O�%�鬗d���M� C�=�v��P�w�b�R�[/N�פ�>�ǽ�0�)��RT��_�t[�Ϗ3���0�?,�D���Ԫ�tKr� 皽���:�*����D�X���b=�$����?r�;~��u{0�0a�n+�x��_e�^�R���d�xFʷ�	�.����h$#��Y��b���A}C�|�^���_u�
�G������)�y�1I��!�.'_� ���)$u�7(cW���$rf&#�s#{�B���Rӊ��{��hY�Q���Y9|�m�~%K��Ǳ�mƌ\j�.�>��YHU�$�{�$��%s�J�P�3���{��ּ���j�{��q��/Y�� �}��apy�����&S&�����M7w���5��^�=3&�(F� k��(�Y�̢ۇ�h�G(��=U��d��$���C#�<q�V�πCǯ���k2�<o�y�4�����s�w�v�(�u�+�}�	�oh��\�GE�ﺜ�@���g=���D}3�Ţ�שּׂ>�g�)�M�����r=5?L"���.������=��א�i�*��LG�Ƕp������Z�-,�l�&���EMנ�ˎF�@c�?G/��S�%f����9����C���4B��0+�	y�;����!�Ȗވi��V}(�FYp>�Ua����&�+��͹��o��w�AB>x�!�e��1����钴xa�p[���7�e���`���	o	�}���R��r?h�S-��l
���Am�)�U�1�u�=^b^�3;ڵ���Eb#(��p5�ϕ#:�;��J�V��������I��>ͣ(fPz�j�	�6��������Bon��'/���@R��9
��D}6�v��X �"�{R�a��KO�@�O�{k�-HC�ҝ�b]�V�<IW�v���3���*©�x���c.҄�--'Ja��wna��}e������ԡ��LϠ��u}���%��O�z&J�t ��E�����@n�F��aM�2I1��f?�mW� ���:ۉ��ųl
���_ �YI��)�����0m��67�����r�?���xU��I1Ҧ�\e��w#)��������V9�o[J)S)�q���&f-�vȠPRŶwR�C	:�8#T�L-]&��z#`���{j�z��_��H�C`�zm| ���B{��+w�|GP!S��`�7�o������tT �0C��w�������\��_
a��I���~�+�!��,�F+�;���)~��k�n)��6|�T�����^��t�r�s�c�%IQ����[�=���zY$k�-�j�-�=�]����g2`�f������#ΒGv
�8���?�񽩫�����Sߚ6A�!�46y?�&���ƭ=�
;5��րD;y��8��|��34�X�=��ػ6۩o��m�,ŤZ�ӧ��@����`�vq��3m���^���D��~�o����_
��R!�7K+ �ɖ�_����rE���?�q�藔��G��=��y�1 ֚��nhb�cU>
�+cǪ��K:����|�@��Ch�dֺsL�Μ�CC�תc�/{?jb^�pa(��\����:2�����hR<Z(�	���J\�V�>���1P=xP� ��;Y�  0y����O�/���>+�.�� ݲp�'t����$�s���us�K����Lso7I�Td����{�\L[����2�H�ii|N�4��3�S%��ë�u,���ÃN	���+Txۙ`5�e-	*2�C�;^��nĨ1��������e�rЊ(\�U�Sbɽ�f*���Ha�j�X���ˌ�^=����b4�e�����"�|�R�N����za�=2g��k�˧H�M��y]�4�'8�����ݫ�h*y=|��o�n��:a�M>cH9���W6 -lv���_��<L�I�Hn��� G=��^��w�%_�Wh���)V[���'"�����v��s�gA�X��يJf�N�E%Ɯ�*r$AA�t�3�$�'HO���W%�2��.
߉�rqGLg�-]W%Bܑ���hdk��;-��g5O���I>��c���R����d�ȋ���H�c(��M� �0�=���dp��u�B~鑽�A�~&Q���E^%w�w*�*<j���wĉ, :��^��y�xB��o�Q����Ȅ{��;&�]?W��[5���,��>0�g-D�0����a�9��ӕ�v�	�f�t�5+�I�b��p?�~,*:��gÞ\7�E:=vrE1<'B�A����i���#�r�K��D��'��W5�k����z-M؉�r�#�|�]�피'�������*��4���1����?bt���0r̄�yq�ʂ^k�.���V\��� �	�u����j<�U��Q�&U���1ĵ�YdP���)zJ��\L�sp\���?�Q�r����^ yP�ݒPG4jƄ;�n�y�.��τ���L���p�R�0h��3��X��<�s���m'��T� *fMޔ뿳3J�KJiBRn�D��y��B��� �<��	�2��dVs�
U~}(~���Hp��bGʂ�*P��2$y����A�q�B4��G�~��h���Ř�o��>�E��Ji�o���.�}v��/��C�K&�4;y�EP�7�x�G�AR�&P���Ҽ��i���%`<ܙ���g�݀�?հ��-��7��V�\�Dػ�6ly&����%�qvxQ*V�{�C��3�M�T��
6��a�!98A�"��=�sB+�����h)!���n�:��eY�{_;O�p�ރ���\����/H�)����Cϫ)�`NV�
���zQ=�:WeJ�C����U�̧���E����D����%���4� :�}���8��ʗ�=�Ū��C�5��p�K�����Ld���$�nEOk0�MfdQ�rXo��:}*T��̿�d2����"s��p������{x���a�}�ٯ�"/b?��`���u��Ȼ�6P��h���ƫ�M����3��/��P��1�@q���*6���u9^�m
e���[\���-��Q��ѯ���4憼.��ze/�HQJ�ʸ��2�A��x�&R�!�@pIe�D^�.IgB  ����%S��0��<Rd�Ռ�p!Q�Z�D�9m���=o��!�o��|-���K�9�F����
 �Ba�	tl�1ʃ+�S�<��D�ܡ�4�EvL��Ǡ�+��K	s�T�ԠL�B(�e}@�ԟ]]X^�I��p��m#	���Nt�f��B��bv&���n�=s�i��&��S�ߠL�Vu��.�uW�b�ܐ����J{��1~�bN������b�b��r@W��!Ee��skYyo�;�6[�(�G-Wrj
�:ˌ:�\jm������R��Sxd�c��:?��%�]�q��bc�^~-���J�{�� ���JMW���:PyG{�x�JE���n�f���OJ���Q�dNw0.?�' n�g�\u|�f�u�JBT���)�!�uz�,�\�8
b��_��$!��V�j6&�"s�g�D(Λ:�e�ͻ��o�o�*���K�_Ȏ�I~$�t%L�b�f�J̎O�"�Oi:�����������2-Q�GV����S�݂y�I�=�t)n����F�ߍ�.9�7n�*�]�9j��ҀsZEA$� �R�zUS�Ÿ��!��7�R�	�`�lR��,7�P?,X�#&���)����-D���F%i0����,�M�2���QO�����x�k#ǝ�y�=,�:�i���V�>�h;�ܮ�����*:Z�3,߷�6�X� f�˗6�#�9"�p-��+��Q��zI���(��:��ڡg(Fx������4P�X�82c�u}\�C�Ъ́{%��<X�R������yV��K���"n�P�Kl\[f�^���%	U�,���D�E�Y��}�weƸ�J�J���� h��QȾ�����g�F��Q���و�vY2S0|����/
�a��k��7r�}�v���O����
<�9�GR�?K��*6�w�u_�;��'���>}m Hɔ����f�)F	�2�n�O�f�!n����5n��ar�-�!T�!f�ZY7{�gW���",�>��$i�\69�6��������A�T+���j��Y+IZcS[����<us�.ן*�3�E{��n����S�Nt�&r�ʄ��6}�1�6��"��SX��	�[��GyEʊ�t�ҟ��1%���2D��kbD�9�N>`n�5%|�-���O��t��+��wZ����<~��cs��r�i�����Ü�JL׹�+hNG#Hj9��:F�QJn�����;?7���[|s�J������(^g�'��,į�V�Ś~K�U.4��2r�K���k�|n����w� �ӳ�a��{����r8�BbGa&.D��`�"��$�"	�!�q�ۇ�la(�{cubZ��#x7���7AѨ��t�bAv=��\�$l�Q��<9�d)�
��`�WEft��E���"�dQ�>�,�'�����f~�hu�Z�7�}��FN���馼g��a�Uh�?������}ݴ��7A/й5aUY�d�%��K��L�2��!��� P��G~ͪ/A�J>�5���r%��QB��o~�.H��X���W���i����#�7#i��2���u�Q��1�&�u�H�{������FMjv�lY��TO����UB�^X���L��N��S0�a;��mȶ���[�a���;_~�'�v���k$Z"K����0C�;)��NIgh�t .��aF4��t���,�����CęM.�����ʱlQ~�'��&SI�� ��i�FJ���ۺ�Í���&�yh�Q�uz���S��� Z_P�~��.��O|�)i�Şu��D��MK
����}�y���Ew�N��{b	,Ē���b����V\QPzZ�#-��?���Fe K;��}�gl�0GZ)����W�W��g�g��T��`Zd�IpN�c�Zi^�>�{i�?=���`.� W��'+|��ҵ�t�&�-ٵ��5Aw�dF��iW�Co�_����i�0�Q=�r*�	��
qΖ����z��-��W�E�粎L�#<�NF��£	]�9*�S����c�
*X|ҙ뿔?����g���ƫ�R�r��蛒�*vk����U�^��Y���Ň։=4H��^4�%=!�Y��4x�Au��n΅mpF���R$��Z���`s�S6<�o3�=I����A�ݱ{yH[UIK,����}���m'?���	Dۛ�؟�M����\�����@t~ޞ��6UF�*�»K:�4kE"�(,�:Db�?	����~��?C#D�uD|�4Pkd"<��UwȾ�sA�'勸�<^�M����A왋��]�J��������z�6+�d}`�:�9��֧��_�_C �<��~ZI���T7��=�d�)������� Xc�?[�\o�o����9d����'m��I���P�����迡���ڦ-o��g�o�8�#�y|��*)8iK��Z��x`�l͙�z�5(/Z���������{�Cdeb�!N:�^@�1v����]������Nd$M�{�'�yB�%0J�0�ӱ�����pƉ��8��R�+[ǀ�X<8�wT�%ɴS�=�D������x�nb]*����9�P7�Z� _�Ʊ�}��r|�O��U.�0$�lmt�n��|�	,���_������6�r��x"��߇E���O%{[i�9��fq�7��a����OLB��a��L����B6_��+AC��O޼�E���Q����e%:����܁�0��!�a�5�\p%gS+�;A�L.B�m�xA	�r�<���'��$����v��7�}�4��75剠m��^�8��j��S[�s��	�d|��~�)�����X䤕����Y���_��	[�|5�-g������̴�r�C���[���(wW�Rj�e�ئ��f���Xϊf�m�r�@�
���*�g�f�k׳�yٻ~g1i�AZ
�����X����wC�Q���K�B��l�뗹I	I���0��� �T�@��؀2Ӥ��K���ꮏ�ۂ��R��/�洚��l�!��bC�2M.��r8�Ex��܄m�9�Ot:Q�P�x��k铬�7�v�eE�';�����)�+e�B�\���Hv�񼕪s���-���2B��ŏ�I����`�&MG�P&:l���IS�1j˭U�G�r�}A��'�W��@Ε���C4��=Z�m,�:�*x��18�ʣ�ݑ�eM����k<96U�����Vl���i�e�x3Q�eF��T�n�H��-w�\���7mW8����/��%tc	$Ed���8�A���0xR��H\�(y5�����h��\�(�a�%�u����>���5).U���w	oo$^�K���C�U���?6t�>s�q���I@y(�� ��$Ϊ L�:���MBNヵd�_9U�Rh�A%�������/BK(+=��Ss��<��La�F�(��+w�4q��b�#�Q�J !�b���P�6��GC'p�]с�SMP�-�����s�D(�,�/d Vnn<"�TNVZOb����َ=��#(,�?H@"�A��k�{�Ŋ:y���P�m��$�Z�����(`K�s�0�o6/�������� +�Ec�"��@dpq;~�|��-�6����)�0�(��&t�fL2��J�%l��L�.-�(�E=���l�%�(���L���kwO����n�j�����M7�#��� ��B9�%/Y�:��7ޮ�f��Æ]"�+{̉')Ke$�T�b�>�[���ٴ1��S��+��R~橆Gv��߃�zP Cҡ	l�A+�h�e�N�0y2K�D���u�1Ꮞ�6����H�*N�J�NݎJ���)�Bg6w���D���Ʃ�,�g��o�L ��%�Z��f_��X'~�W� ���l���5@���D_Ϝ�DY��偿��~WO�Y�p��d�����!�5�_��h���?�,PI�w�enU�f⑟�v��L�2sb�~�2�
���MdF��׋�P�%Oh�E�s��馿�M�ˁ8�dF[�ڳM勠'ʢ�ttf"����>�c��e�ri�!������ok�Æ�o��,)7Y�0���2�h��C��+�;1�uK��F�g�%���m�T-��� 9�`��$c�B|4R~4�.MlW��4�+	�ԣn�J�m �ۇ:�d����Le��
����,g�`t�������� o���E�bX%�!�μD��j�2۽ê�j���8���K	�`��>/��ُ��
(�����k��v6���r�����ʹ�U�[�z;jgC���$_��<�&a�y��eA�ף�HW��[>��(���J|�X��Ě_?,{���B�"�q��@G�}iL�rk�$>"���˿HZ�LMW�~C��m��S�Ӭ��x��w� ��7}�J}ʛ�����' ��C��C�~m��yV�8<e��n��ܺT��cf[t�Urv��؉;v"m!Z�9ە��ç07y��	3,rg����z;9Ў��|��w|-04�O��'��8��@m��Q�06gUC2���VE`Kn �ctB�]���Z_86?��÷��|U�{Ԇ�6�[suw>E�x�~1���m'xI�_������c~�'�Ѩ�z�\�{�+g���fq����߸�_Z�u%F����������\�>秮誃_K$��פ"h�����``�>�Wx���Oi��v���T*U�Zv��̙���ﺁ�|3bb֟��(+����WI�{���T'�=f�\���=29��BP��)g��Z�'jJ����8Yk �D������'y�k�{�l�n�v��'f��M/����j@ڱR���-����<ٶR����&p��	�m���p���	�l�����)*d�؀V�
���Q0���Z h�~�D�����땒���G�1�4ƚ�&�ŗk��f���ٸ�ӵr�ⳁ�3 ����ɔ��ŗ����D�5E��o�t��ȉ-����6�R�@=���nG��K��Ht/kX��c�'�bz]u0x����9��X���ԭ{�����O�9���zYQ>�%�J�u�2�FEO�֟q�U�+�w���ĭ�Xk�k+)��3�wO�W�%%2�9#�_��}b0�ܹ��uߩH>�͎SB�Ae�/>C�rer�9Rb�B��ʀ�	���F>�l�+g�q�Zcc(<]ˉ���ǜ��D�l���'|��G�_b��7�/���r��c�b����+-`#���w��b�_�rLi@5�˘ A���ۼ��J@cY��#���'���3B����R��� �V�թ��s-���OA�J��K�`��!_,>jO ���s뚪�Q�~�Z���W�|��T*@���2��
P���ʕ���x����x��ܵ'����q��>�FlY�M���ݓ�^����Ƿ=%3N!N���H�;S��e'\h��;J�4����v�E��u�`�9�x�tcM�^�s� J"{��`<��h#�6߽]	���9I�s�HD���h�b5Q���=lϿ�|?�]�aR9��_�]s���S\O[`y�L� ��-�&y/I2��B�ٲ��ܰ��)�(u�4^��P���[P��J>J��-��c�����𴆛	+�ɗ�d�����'��|U�o��a?NK�u�hc[��B'�n�υ�Q�C�,�1��Y&�Od`̮j�������>f�I��}�2/���Ww�I[�1ꇓZ`��S*#�pU���&�#I�$M�Xk4�0O;"ٖTH�D�(��0�|3tEB�9�ݎP�v�`�w��;Y���>Jf�R�S��]��Mtz�q{�k�J���Zl��Ί^�Яa��@&7��ݴ���.b�~��~���E	���y�þ;9��Ȁ?<p����ʆ�?�S��V������냘-�3����虹&���Q9;:Ӻrc�]�ﰏ���cV��˗�Z��&�=R.D�ŋ�(�v�@c���F2/5D�.P+S+l"�.x;V}���t3�d^P;���p�A�{7C� �r�1�A�5�!qkϞ �t�C`d�����g��櫌�����,��K�\�V���$�?���7L�CT��K�����{*���9rh�� �֞�������¼�}�I@�w�Z�g���s��T�7�T�x^��s;�<T�<`�=��?B�W��n}\"��N���c��������rʟ 9`q�6���ܖ��ߺ;_�b��&���o[�.�A�ũ2�`�v�I���WC2�
�x�)�XJ�T�(G�^�B`�D�or��끡���Q/L@�w
bٔMI��6��(�7g����ˎ��yMb���� ��7�4���@u}� ����ҍŧ-����v�ڈK�0��'gW�ҝ�jIj�54�k��з9��P�A\�t��P��|T\=h�-Nm�p����+C��K����? �����01�� �*����A�i�U�EW�T*$ G��_���-r،������V�+X[��jy�*�8�s0K��k盗]��QA��S��g��1�h.�-����!Xf<�$�E9	ϖ�g~v�o93�n+��&�V�RC� �&�M��(�FL���8���E�'�ecdf1�M¤�.���4x꛻YTO+u�ZZw� �g��=y,T.#vg��������3�Jݒ�R���[�m8�$�d.���e`U��n�R���C�*��͇�K��5��W�tٴ�	��]��J�6������Y��J�0��:Eq��`@A�b%'zO?���4/�ؔt�rq��\��y|F�rqwa �?m�W��Xn��=o6�ݾ�ځ�Ķ'�;9��r���?a,x�!�C��"]=���bΗ�Gң~���O�%|޹�ZZEV���T�EQ=���,�$�),W���z$�5�;�l����t-HPW{�l0���C��O��3���Dv��SLM���uh½b����JY�=�,�� ��]8��@t��*�ȗ�2�s�F`���I�<�g-�y�^��?����5_�$�6��N��̌�7k�"S<�/X�q}�x�l̃��.�=����T�N�邗� ~O��C�M����E�r|7�.�� �X�ݷ�W�J����X��;�v�PE�{9����W�i�r���䜙`�9�hK�>z�7�[91�K�!xg�=GV^2������2q�����tK��Ե��$yw.���K<ڸ�X����9~�^����h_��`�4r�,�P�F!&)�*���g��ӆ��X��:�h-Mm�1^�"M3����Ekf���y�h�@(���U=g�x�U��Ss\�����3ϧ�J�*�H;Z_���q��ra��B)��c �Z���[��V�r �(�-ަ�dȨ9)���	�>�Yt��V����u�|�]����!{]0g<��$ꖦ!�<�"=����ۈ��-.GablYx\�������ҁy�I)�
���Zع�M���� ���S�b��_�]����@��&�P�N��Y�hk<U�O��z�饰�f ���=��P�;�}�ES@�ſ��"�,=�~<�$1|������s@�	�6jD��(>��)�6�B�@n�,�mC�������kX�YpX"݊#�ˍ�w>����0���C��%z�c�l,R��e�Q?��(��B�1ƺ&rS.�~��{�s>9������a{���p�%�S��F�ʓ(��߂
c*��h/T�խ���@�� �;� r#a��A+o,3;C��Q�6z�����(���>T�fiCڊ����e`�!�^ s�s�wׯ��'���M���VE��p�
�=sb�?����r�����}�.,c~��K�n�;���f��S*��@v;l�����Sl����|!���l�R�J�4?��۠eѵ{+��7�,6%( ��bi�� _o�c!q�&/�ͮ�z�ݷˡn�	�Ϲ�z�#�_�9&Z�K܉NC���ِ���u�KȺ:�#Ѓ�G��ݻk�P�l�
��b����;b"0VAOO����L��.�@iܼ���֑�G����k��	&T�`�>޳iw���AWA�����w���5�hl�hln�[���=L'��M�Z��Ԝ_�0����e�E"Zi�U���;�o�@f�}"m��>$�R�*��I�_+�K��jN�H�ԝv#�:ݡ��m�Ʊ��>��gR��o@<$�7��+���v��E)s}�;59xht0����e�3�~8����.`}%�P��ց��O�l�����
N��o1MJ0��Dr�Q��՞�?��J��c�1q��}0��T�,[bq�-��,��. �J����!ĵB]Ñ!��FI��,t/�񬮓vS���a���-�x�&�1ZU��")Sǀ�Ӱj��Eh���ڍ�й������
�U��Db��?03۴�%��.ki�N�Y���#��J|ޓ[6����vJ3�b�pӦ%֧�X�Y=����k>��u��Μ��>��I�`�Ԣ���V9#��)�I%����/%���zfRi�߀������*�fF:A!ks�,Ec�?T_j�~lV��x#�T�W����U����W+��U� 9G(lľ��k�D���9�z}��
�D^4�J^h�}.�����
2�w�\Ӭm�hkY?�G5t��_J�m�-2��H��-��)\�e��f�S��;�+�l��Bl��?n_����gٷS������ ��|n�l��wX���]��O�H	�(l�oIZ�?�-�Mq3�G�{��=�=o|{��0�|�MU�i{W�laef�]���m��v��%���X��g�7S[�b��5 �{=*�Q���
�������%0\џ_�l�{�Z��ƪx�DC�6tڠ���~೷�hW��i�F҇K*<Ȩ�W��^�	9��v�� �3����]�U?t�y�E������m[�}�jK�i���~��!c�E�0
��\�٭�x�ٛ� ��05-�;̙�}1�H]_��	��>,�貣)����z޼���I<�eB}��1%o@e\�_ZI�IY�$U5��{Xa�o��<��cg �8ɈF�Tc5˂�.�Sk��t#�}]I���	9?t��!��/�"��?I�ڏop"���6u��i��8"i�p�������3̓m���q�\��{cUᒤބ��R�y�>׿�>�g�wݠ&�%NE>	�=��o������^�y`i?<�o��qp����>\�o��R��?=��]�5�^g	�|�n���� �
¾E�k��4z��H�홎�M�H�Ghu(�O�� l���������ҧ�Fm�q�ŚpՋ�z*~$��p[�R,�H�ظ��}�0s�).q��/�h�J "��b*�ք�|f�x�����7�m���ּ�*J�55�~��vJ	�<�#\�6h$��#1���bo���I��ʱ��C�t�pV��Af�o�I+3.�bBk�����eZ
�F����t
��o�����o�B����@}�_��}��e����E������6B�+ovvz�e���:�a�ұ���M�ɑ�E��y�`��o٪$���jX�e	���z��`���b�>�����@�Ac��`x����*��g��shUIMG'
�����K��.x�׳u�����ِ\����*��:{2���v�E[b�eS��̾X���o�I�&BC��g�䮑�^�:��"�~~��S���뾍霼c����ʙ�l���$x������0FtH(Ѽ��]�|�r%CZ�~||mۢͰQj9��?.��<��l�)��)3�2��s/T�U~�ж����(Q|�����	Q�ϸ��Y�������V�Կ������V,���+Db��o	�0b\��i� �f�$��8~�6i�a��\��=2�B�����W-�F��3�T]�L�N�v�H{��{�����=������(l7�z��3դ�@R��C�u�`���!�zY��H�1�Ј����4Ҋ!y�]���e=A�����jS�D�w�4d{]�����gH,�M�SX�gs���:�W$7�o�fs���a4�w��m��!���'x��s���dͽ��0oXz�M�+��
��Gf	]3�#m�9��bߕY�͜s�P��2�i���d"E�2�g�G���_/�CM�u�� ��L���=Zn�l��.gEew�TPE'_!�S���Δ΁��@( ����Z��ؐ0չ�A����bS��$��3����*J�Ƿ��KW�l��f�Wh�u�Z��A�M�1k�E/NS��4�4����'xT�h)�Tmn/�@�Q��U$��tJ����hF���^l����W�s ���ɡt1;��]�t�Ku�����~x�㴽7`'Ǹ�Qx�w@�|ZZ+ �,p��4a�Ƹ��!o�����,��| 	P�r�]ſ�9�e����z��8�.�1}7���Cͳ�2 ��b��?*P���Q���O����X8�~$�I����8-�t����Sp^��f_����~p�x��P���SC�ѐ���Ηʌ�x��}T���"��ON�iB����¡����޶�����/Z$��U�θr��x�K���G4,uH�������Z���IhxFC$6kq��&��� �M��eu+o0?�5���Q������Y)g,���܎��(b�	,b6ue��	����iw��7CF��A�S}.��AJ�Hw#�5���B������&�%�	B|#S#v/��縿�c �ohq���-:}�8V��O�x�{��-}t����Z���{H�4�K�o/D:����Jc���]G�CU�A�3��V�DGδ�d�9rܳ,��K�s��΅:LMY҂��_c���Q����_~`d�������EsT��G�rnoP��t,��樨�]-Vzd�k�Z"�f�bZ�ԴKƲ�Qe�f�֭���]iw��q�!چ����=�~l�É9����>�W�Q�4ԍb�����[[�"m��UZ<��������Q����~a��_'�B�H�J};:�7�z�R�b�$.�����W�@&��vXԠ�Ru?b�C�x�)�J�b�\���ƥ���A���´u�k����������F��-&�������*y�����(Szp�I7���n���siM�_�u�� ��.�0b0)�σ��_)(�i�Oem.��b��>g�KFb�/F��/���y������ʫs�_�Ɖ}"��{VM��$�.�{�i��p~��M#��?���҉-��y��J�F���2N�P=p��@�����U�vHl턍d���ˍES��EX+����ݪ���y5)��+�kp����ԧ�mU��������T9�ȭ���aU�>EV�L�!���DtKo���4�W
>�w�:>o e=���Z<_��ѭ��'�]Ɂw[߿l�@��~S��Z e3�Q.b�{��n�,�I��,�0	��#@~7�c¦�������GLˤ�牢\��Rʏ�~6�cO��d�EPV"���3�aN��R��s�&�]� �	��)�Q�*�ԇ�u�O"te��"�c�f���>��Q�.&��_虜��n�a��!::��׹
�)�� �#�EM�$���i������EA7W�|��6�<s���CrRQ�S1bE&����{�馍>��Q]�0x�BJ�j����Ju��}Ml�~���W���f�r�9u�hbC�`y�!��'9�т&v�X�a��C@�`�� �)0}���$k��z���]7��Z��~�~���Z@�=\	6^�F$��ґYv��S����T)Me~M]7	:]m#h=��50�2o��Г�pɩ,z^����`���%l���$2@������N�ERsm�C�$NeL��}�.������	��dX�=ئ6	;Q��J���Rd��#  ���X]�_o�E�c0� l_[dQ7�>^?��(%4�ԕ-�H�d<�,�{zg���4Wy��&����ۡ��nNȟ����t�y�T�ϐ���{�{�
p�V�1>�0�?]y�$J=FL(��q�J��J�p�@=�=�R�M�f�,�ٻNb:��p%2G�4xZv���䯉de�P��i)D!��P�m!�Ј4v�ﱟ�ID�Bx��XX�ԏ����@���f|�c�D[eb97��.V�T��DCӺ
"�dN�/����h�i�'�N�hك#uS�C	�s��� oq ��qX0Y���Q[���*��N�qP�W�=Rä�砥	�ÀR����E��{��Ne�c���g�s���nH�@������M�������>�E,� F�	�"0�NXX'<���n]��T��Pv
S
D��DU��5`wq����g%���8Zs��$k٣��xc�7�1��t�C��j	�G�K�&�:/r�BT����bԮz-b>�V:7��^v
ζ<̵M��G=*L�'�)���FaY������uK�r"�cV�����o)j#�+�N���|��,$���+8�:N�}�������4���:Ŧ~8E����Ev^�I�w>(@ME3G)��*���=#K� ?,���j&�^�qG�;5OB�21>�a�#:{Qؐ����� "�V�\�+�� ���D�����=�1�B��/���C���GK}�J��5`���=��_�L��(���a��N�,&���h��>�6wm���J;B�;�m�A���
�"�s�ЃRˍ�n��Lq�3Ă�	p�e�@�F��dOf�1�u�R��(��
گ����{Cz��q��s�R��d���8�ݮ�"�n.���"�\ E��	j�B�AҌnz֊:W���Jy��{�1���A4&/��c6��C�X� �a�}l���θ]����u?��ҕL�$Kh��z����qRi�:�[���/H"6 �D*�蟧�pߋ�4љ���
�-͆`r��w�ts�"�d�βRHTJ�8�-�N��}��a�V�Qo$K��E��Jy�E��xtq�GOl��1`���٨��e�FPԡ��!YS�r��y�'����?X���&˲J<m��|�#��jtc��3����Z���WT��G��w?̩���˗H�Q�+d�I�Q�����ؓ@X{���l����y��C`"��R�vL:�)k�?���:��&�Yk�q�b�:�����3k��ɳ��OrO��T9��@x�䰣��5&�h���(�_������iʶ����Z��<K���ڍ�Z��>jq��i��D���'�$%�s�z��1�C7=�W[����ʗp��b��X�c�ڐB�F�+4��,��s_�K}Bpyq]��D��}s W�q�x�$�񵹾��-a� �r��[-�.TSA3���Z<�.�&k;OIo�����=ܾ���%��}L����K8�"LHQs5\�e7��\"�}2�ygQ�w:X�M���W7+�lkl�i��M��ۃzrG��Y��@�`H�o����{|��:u
{���!�O�2�0�-G�7/_-��`�.k��Q��'n��)�h7Em3D��wq)��09�>��q��7��ơ��#0Z3�f5��=;ON�6�{32��&�.)4��1Z�-�>�eK$np�ʿ��f��u��&u:$%}��.hi{W�@���D� ��3�,Y�A�!��C@�s �'Y�8�Ϣ�0���O�2��،A��>�-����N��e�{�E��@�����S�qC�8�3eT�OC�I����
;�R8u��n��v����߆����O�<�ʇqoQ�c$:ki�YP��jD�c'�Q�;a�C]n�7��@`ŉ�	�}2o
�ҚHp� ���lE�����`��)�Ö(Z��;pO0��G���a��{�y�\��ϺK�ғ����o���Ӑ8-�oZ��F��݃ٷy�s��������&��?_6P��G@A;��WJ�b�*R����X���Ec���F|�x����.z�^g�����rM���VD��]|��aC ��aT�m��ve�|חa���1wI�I�����><��*b˥�>�̃B��P}U�b��ݮz�M\	7�ndCC�p��ڸ�[02V+d'�??��}�R�K���Q�I}u\2��H2*yhj�� �T� P�3H0P�%9�R���;r� EC-�O�z�Y�"��Q�R�貀$-_Y ���IeXe]K?�Ҭ�M��$ӌ�@�'Q�9���FVPT)'x�Vj��˲Y x��9ˇG��Df׳�_��-�'��_��Gۓ��}���]'�Ёj�������@�gP��6ԃ��� E�q��D�e�.��\:.��
�s.��׹gv8�i�Є3k���o���n++y=mo<���3P�y�ﻣ���6��<��+���d��-k���(��M�q*�-�1��t�*c�]O������ffŝh �f�B������b�v�Q��ZN�<(�|}>Z��ː$���7��0�m�m�:���5�'�
y�%ZQ�(؀A&$e "�Gm#���w�i�8�qO&���' �]<ڃp1��$|n�k�y���Z吰>�E�o��!Y�����!Rz���#���L5�T)�2�&���x����Ǐ>�4�Ǝ�|6�+���zʂ�]&�j��x�s>�0�P�n�6�](ӓ���v�ꢤ����n\��Є��H	0�ǖ�FM��%�u�N�]v+���J����=���%d��\dGEh�UMN�Sv�z�������U,�4d��P�M��dy�Ó�W1! �R)�F����)=`��e_�N�0��0[��a>CGC�dQLnv})*�Q(W���� /hSA~}Ȝ/6�Xi����8��e�����#Cj��d�:��en)DG5��D_wx��(uۍWBpuPâǽYw�:�?OM��\�:�<ܣD�����G� !��/𛲏3F�5�B@R�$O�&\�Td��r�ʏ=�8� ���ܝ��!mA���[]Ge~���d?Dk�����[(�|z7�ͲEi}i�4S@3����Nb��*8�"�/k���,UH�uT��ӣ�ov��{��s��WM���=h�N{桅S��h�t��7c(/��;��i]$QU���0����v��j�+?�4��\�������$��44*#ap��\���Msc��qb�;����م7t������5:s��{�����g:�f7��<KG�e"as�6�Nv	e�}��;9W�J�[�p6�v�ݭ��9�u�8��7	c~c�^���T���u��[Q|��+�߹<�cZ�k�DmBȺ�v��M�gC�)���p|>>Hw!�V����h;��$dDs���ڻ��'F����vcf�C�F�4#��}	�6_ʀX���9hj��nyi0���7x9�=�|��|-EQ��,�<�:�H#��K��+;��3$������h���@D�<���&�����j�=!?x�}0H��;� uP�^��<�O�9�Si+n;���AUX}^��҃=��ǭ�\۷���t���t5���Oh|�?%%��P/�ǓƉ��%U��ǘ�3q�ǬH��ycʴ��h����F�a��$����kǏYUڴ�t�3�$H����ͮ����P�u�}U f����b62==�;n'g���3��Z/�B��܂�$���Lb�6��C�}[�㖷i$�jvM�*�_��%�֊b�hf2�Մ)�r��&�V�,q���s��%�ՠ��C�9�,w<�o���Z��O���Nh�Gg}��Y�@9#؊	���`f^epW&hݑRP�ϴ��������
�Q�{�~{�kT��ԋ�O١)��(33t[l�fl�XUl&ƯҲ_g��	(��z��b�X��	�a��mó}�3�gz[��PQ�4����g%o�b[֔�%�Y'���:���Y�9Vx�V\	X�0�?�M�c	� E���}C~��M�h�G��5o�Ş�ֿ2���ڡ�W���m�W>�I"eJ���1�PC�x�Fe�J�H�>>�6��2[��R��ig�5jŹ�ɮ:���������yˬg�y�W�Vi~�^�'v����|��L�K#�ę/g	��y�5t#��bc����,��U�� �W	wCؘ4�	�πե�h?������ȧ'�� 練$ ���C���K��@��������)�6>H��J���C��)�	t�09��3<�p5"Ul�ݴ7������v�$��*�밚U�p&]a������F�+�HZ�,[����d����|)��UM#%���ӄ@��V�lm��D���
��.+�hx�X>�Nl���@D ���r1��n���[��A*�����ODzv�Q��/��	�6��ĤK<T�w������}�PAGL��i�g��Y��s�/z:��
�E���#S�� Ʌ-m�~9`#��wTO�&���0}�m��R���/�+i�Ê���R�[q���Yy{��~C���d���t���7��u�Ȃ��,�o�6T\�Z{�U\X�|=<³k����Qשc�ϋ�z��,�l�E�Q��/y"�|�\x�5WGh%���,��Uc�'AG�������w�>�U�;G"d8j�SNm����t;����WUs˨Y�]��<�� �{ׄ���3�N��8��_�'v[�V+ml P�����D�Z�Cl�����e&�:̴����f_�����*��m��)%VF��>�\��4v�~���_����;�&�l!�+|i�H2�p��y>�K�Y�[6nD���/���bw��g˖I����ꯗ� M%W��J=Z`�h+]GI��ROZ�X�` �o� Q�	�c���g�g5��$�ژ�E�4���{�K}KA̸����%;ך��`W�p�|� N��&zg�؈5�)%T��ȳ�틴}�AEXۜ�-l�� �|�K��70%�j��~�-�}u���ʉ���9�¯���n`�2��hQ���e�Y(����bC�3�y�p���̤�x�h�s���s�έ�0�DE�a��'��0�U�6]Ǧ�n�x׊O�[�����{�/���2@�:�ك	��T�#,dQ� 3�[���|�� �"<0��B�oT#��|[�f5��F�>��r����S&~»A�c��o �k��v-@����f>�5�?S����x.:�;�&���mFb��f�[ScƄ���L]a	�}�|BS�M�F�u�WY7ЄE�ٶ�Sx�ּ�2,���.��G��.���<�:� �:$�]�c��E�TzA��s'�)u&N���������gl�M>
�g�@ռ��J��k��X5{���u�L�-�;Z�_�d���b��+Eֈ^����qū0�B��j�Dτ�~�-"�`�34��B鶗��P���n�քM�sʸ�m^e�.�b�XT��E~������Q�@Nl0�\2�a��b�20��s<4T|iע{�C�a���.���V�8�5��߮�9�&�t�DJ�M[ʰ�u��rX���4-v��3F2tS�� �o�@Է�Ɩ��iA�[���D��$��>��;�����J:���Ï!������sI���M���u�� �������RXTR3I�.����L퀍X����Z�pB��D�V�Z��j�OR���*����ȘY۴)��`){WMo`��0œ�H� �̛��r�m�'�>���i�#c�\E�`v8�}�Ou��椲�t��&m.7�D�Z*���q�=[ÇS�7� �1�٬*?�Q��D]�H���;�9Ԏ���7b"S`y�g�o��#s
�AX�yW��X`� �1.'uӬۼ��dj#'�]+��������N�]�S��7��p(��(<1�}����v���P	ϊ�� ��B������X�`xU�Z�c��8][3��&�����"�[����[�z�̣-�M N��rX��E���sDtv�)��!V�P��	������x	Ĕ���,J-"hu�ƙ\,���JdA!䊓oO��uEq'�N��3]ѕ�rDxfMlG����9$���~�Kϭ:��rߵZ���dU\.��+���Ł{�*�}�E��)��Y��zac���$T$�P>'"���c<m ����Z��"���'x
�2u����d3%;��H�r�I������sB��9q�R�����!�� �N�A']�|V���0g���Ʀ�� j�H��hg��.tR���?��.�6{��%���A��v�\�DNVm������DX�?���mv�2�<D�~�2y��J'�i"��<l�C"+b�n� O�>z�8 4#�3�y�3TS�0`�Yf����4ʀ�p����$*��|�o��uް(��)!����Q��!��^&J�7v����+��[W���NC�SI3Y�-�|��0mC>������uI�:��@={l�%�o�nv�9qI��f։O��%�|��$��{~� �J����1x�p�^������]1w.4�r�׮&��n�,�cYP�k�e� �ή#O۩�%z��ëjF�U�C�G.��V��6�>�5�a��%$�2-��5��+J]p�tΪ(�����]|��qGcu��Z�U:��ύ�X�|���E��y(i2�6x�{?��ѯ���fK{ZN/W���Ud���TO�~. ����m�'�A���f�$s~CGuOi���3�Y�����X�p�����;a/f���U�nu̦@%��X��O&yդcr��fb
皋ǜ<p �?O�2݀#�B1�Qq��s��w�g'+��<BG4OC[�^<`@���D(dVaaе�}at���l)����~7��DO��'
[�~�"C����̀mZ�����H[����P7e{�F���(t#e5�M�ɢ�}K�N���@��qxs���z�=��u��T�_��b� �I�T���N�S-�V���l[v�T�_�1�e:Jp����h�����(3���Z=6�Q��E�������� �6�����`�ɭ��咽*���,�1��]*0͍���!)��� ��1 �)V�*���Ǧ����;~��#�����z>���U 4�A������%y��Gֵ�07�K\�v�y�󳚒r-t)������ͺ��~�!�V��BN��f	��^�U���<x�n�BO��_��;��o�M|�8&X��J�Ĵ�ܷ�N'ń�0��@4{"����J5x�֬r�0s��������%�0�|쇄�݅0V�z�$�k�����\9y�fThGhϢ����e ��M�G�Rky�,*+�9 5kΔ�����#A��Q�_��7O�5n�Ȏ�9/�����|���G������Q�,�Q���Y �s�vyc%W�yw��/[�|�� ��c�"H�.Ɍ9�H���vLL:�N�F�w�Z+:�8�HQ|��A��f�YײX����c�8^�I�8��N�*��S��5N���|U�:�S����R��4wl(����(��
eh�?
�B�E ����0�Y!�L�( �^۟����Y�F��<ζ͠�)@�dl����X~�ܩ���V��g��v��j���b26Xץ�Vk��XنrN����qO��@j�b�n��G��<��\ืp�N��>eĜl���Eܤ����4My�o�\?����VfMmٞ?�CЮ��B�,��'�ߵ���
2;t��v���르�w�D���e�鎰z�&�!S�M(�xU���n�/J�������<'�$3�,u��w��̹ܼ	�� r���y-!�߱��f�ln����V��{�7����}��-���4+ֶ�:���~��x���+�1�Tnc�ʣ���4�6θ�&Psi��Xe���V<��B�u�p���C
3T��z�tٌ1V���ϐ���~m}4�A���.AE�'`ZT9�d<1U�/;b�l�m�0!�3��H�!�b�q��?1���z ���"Ӆ�M�R	F\Y�����S�Ah�����0�1�C dR����NNc(�lY��#O`at ��"��rlB��
�X�θ���8��
ͷ��ɕ�O�綇�&��;r�Oh�Ȥި)��i��!���?�����k��V������?U%&�ժgz��óti�!6lvhH���53n����n��3z �=�IE7;Ɣ�.�h�V�?��K���z�b)��b�&7�C��&�8���_��Hܘ@g�,g@�taE5N�x�%g�y�������C�Z��l��M�y�#J�:�
��̲���@5�S�T��n�"�w
���n\`��`'$�)S��6
Z~��>X�X\Ρa[�6YQO�:)V�Q*j98\.v�18����-�fr���\���R�� DA��ccyd��2�4�Yi�`c��4e��義���2��7�4�BD�K's�^�ae��3��I�9���˭��}���X ��E�1��H�%��u�u�E'Q��,�O�?��7��p��Ve?4��h#��s%�����j�;��Z ��9��WCI,�i���������̩�u� nED[��^��;��]�D1�~A�����}�U0�&vc����j��wd��ԥV�&&vu��\�>��Y#���#!1g�y�Y0���=øyZ��JwZ�ViЭ�e�`���XEAE�k��*D@.�>�Wu%��|�i�7��?Jpx��}"�.�=
�Q��T���K��l�+]L	�2a���5\���]?
\��%�l��X:7K[��͝�x�������-�g@]x��I�m�2�?B$�D��C�Q���R�%aӖ�OM@x��$�\�JM؆Q3Cm�Zg���~�`	���y�tԁ�]c
妿,F�Uw�h��A�)���@+ȸ�/-�+�,͚l��_`��.h��֯kԦ{��1�i������J�>�����Xn�2 ���i[���f�U5y3	s�E�����
0 ���F�j�H��-?��߳����V�9Bɶm�4�3Pl�b��	S�A�o��.W�~�^�:h�}�ϲa��v����Ύ��<P��'�0rET�kt������L6(i$�Cތ�SYr6Exۢ�2i�?����lx��<�\\ue��o>�Uz����b�7����p�kI��Y�F��R���>�;��?�6�}o��?JUhE�(�-.|�bCc̑�p8�������2��*���>�99ؙ�� Jeγ���7�q�(��5�\�7�J�A��#��/�S �=���)^Zr�^�yq�5|�.�VZKvW@�;�Zg�F=��BaXY����_l1�>�u��W4�|�ڞ'܁Gdp����f�4?��NN򥉟��/**�Sȱ�� <��H��"G�:�*ٿ�����4`�ٴ�v��ᘉ�'"�\W�HPj�<����1�*�b���ªw�@k@�e./lj��aS�D}?*��I��e�v�
���W=l��(���5y�?��]���x	�`G��� �7L�����Z��Q��d���C)�ȵ"���}֖#� �3'-�Y]^���2����e�5����:u���r͚�-#A����j�`.��*��b{�s��6����@�)P�!�J<tw��Եg�[�!�����#�><"�Z��'��Z�8���Vm�jR�eO��+j�뼲���p6)�O���l�������_җ*�l�����aN�,�3f��xxn,�~߅,1��ĔWM��i�+�_�gI2��lˑ���ܙ�б�Mi5���k3�k����`m�&΄ի�H�G����pi�W��x��,r~�1m� pK�S&ݑ��&�T�'y�2���=���c�X;K\����q\��Q4�]hI����uM��;H:�f�c��sҌ�ل<(w��w|!�#���3"��lh3c�!ņ0p5	���X�����m�n�'��
8:b�����IZ�YmѓY��:�}���E�4�n��N���g	�3�n�*$��na���@$�H��+@��Ev'S_ R�	 �,���e(�7DOsdqEţ��5w�V��_�F�e��������("E�!<ߏ���Zk9j��29g�������&-���ow�V��G�&�\�͏��@���;������tJ���O��3#,!�-��cùk���P�Q5Po��ؖ3�c1]F�ޢ1\�b��c����I賡�z:}8ځ�3 ����z.����h�A?�M�� X&�o�������� a�ԭ��֍T�Ij?г3c��){��i�9���2�$���]J�HQ9
)7T\�ߝ(�o�T������H��GF������%�/��������L��@�w������M�T���uNF'z�<��һ�'G _:V^I�eZ���QM���s�٤�,*ఄƺ��d�GY�k�nZ�w�
4J+��'�Ή.(s���"��]�(%$Ҳ�;v Š�!�X��a��x��L=\[�|̯�)�d����TZ����Th�s��DbP��,��2^��g	y�n���j����(��>��9�R�}[�b:�Z���C-��?�A����j�پخ�1!z���=+���(]���q�}�yF�2j@~��/Bv�p_�'a���
2��Yb����::�	$����sv�fw0��)}���;�3Y=W�NS@�ͤLݘ���MW���ar�8��~6',��ɖ]�5�)�ҙ��ZS϶^����0�<���L����ZQ���4��� 4.�\�H1h���
�(0�L�Eom}^3u��S5!|��Y-CC�5H{s������d�ʲ��?$�qlKz_Y�4�o@��Cv�d�Jr,��e��n�>3c�e�����wz�C��7��龇�*���G�CO�k�aSA{�TZ�:*��&����eA-@1�����rI�Ě��"x��ʔ	��I=���y~�{�ԛ_�C��2���KrϮ�wc�;�e*s?
���G̰��q����E_��X�����b5�S���lw 5�ҹȯRI���*ҏ~T�Krr���˝�B�]3�~D]�	)�R�<ƺL�*1\!S U�-���G�
Ӡ��{ɕ���Ac��t���)��8����!�к%//������(k�@Q-ڔ��S�D��9��Ƞ�d�����iX���L���;�VDI!��\T�����	7�'�ʱ0B[�$uH��`�.���0��*��ȻyOJ�F�S}@��y;a�b�����[��C]g���Vb�	zu��b_-0�8a��-Yqo�L`�η#����-��rqG*�s�W��jyF�G]\Z�p�JC��f�%
��ʖun��f>`gG�8���I�݈w�?�%?<c��KOw��p�[I�?������#��t�~7�Pn"��?6┭�<��!�,A���#�i�/�u�,(�k��m��7<��VXF�F9�m�[���7�]�s@���_��5léOD��R�M�7DܨBnER�3��y�n�:g`�_K��X�m���SxW���ZA8�����{WJ+�D
=���N�-�2�G��9G�Ns\�7K|�r_\��̶QL�}_\iĴg�#T������"<�H-ǲ߃'�ܗ�H�� Y8�Z=��ʠw}�}j�0�L侵�8G�� �����*xi��u &?
�+�;����!I�WW��M�&SM�$�������E���и����"^��W'F��#d����K�b�A�D������[������s%�N�?�� �<���]4�xf*����l[��mŎ���Q�,��@r��*���c�dw3��ͅ��S�W���ք���>2�T� �7XT{,\霺k�.�}�A�d�8R��1F���&8�oX]Qi��ǐ\�!���t#6�/#����d���lCC��$,Z�g�o�L\�w��>L�5(�j����g�~R�f{�/����P����A}jek��)7����WQ�ڎ�j����(�}��N�D�p@tj��&��f�ʍ5�3�jŦ*�+\y����/?��fT�$I�?�sB��_/�˼D��A}��69ǃ�=*s��^&��wz��$���h��ߛ��(�鯇.
3����Gh���
�]�����#�%�UO�L7�yy�P7S��M"���������]�F�¼�=��"�\"Z�wYogyuy�11a�!A��Y~�����g{<j+Xa����On
��Ų�s濞���Z�&4� �PopalU#�K�Kў���`�6��ru��n��i���w��_h�sb��wl��o`�kk�Q��.IJ���q���:��l`Q��J%Y0) �܀����R\b�a^�hz�k���"��b󖦃9Tx��y��^9�&����6���iM5\v܀�ls;�c�����'�|~+��Md&9 ��?�XJ�*�ݶN$���;��7������&9p�5�k�ҩ�
���ܕ��C���z~w:X�;�G]ܓp>[��d��F���]��$�̩��!�
C�j{�{�v��x�Y"���w���!�|�~S��?Y�������[��U����q!9�Z�X���+F��D��q��̃�
F�P2/�crDs�b5d��tB'�x�7��O�6?4�/�9],%q��e�Re��r�aE����:��A�d1�'�&^ZP����	m��]����7^�WE�f���AP�G-@J�i�� ٍ#�"��¾k�)�g� �)1l?\' i7ոnQ�o��:��A?j?�:�PHc�MSED*1��E���ޮ��|��o���a���������8ǁ��|�����K��-�r�rL�����۪�?�	�%�t2؝M�Jm:��PB^��L���Zws?��pB�D3p�s�B%x|��
�?\:���;!��L�@����2���_?J�@|t�T�������$��co>M� �ڵ~;��#�Tx^Q(3�4_�M�_U�����:�|&� �Y�<G]�n�q+�ZdMg5�Q;�L7��j�d�ִ�·�\���a�{��js��$�Ua�{��s3šU��?���?9�[�m
&��R�?�9��#�������T�����9.f�z_�ᨋ���&'L".�c�>7��)J��fȺ�{����*��3���̖�*-yyH��t�A�^��x�C�GEx���6�!�UН��`��*��*m1+x��<<��K��L5��gom~@TY�c��e��q>���NQ��l!L�D|`�֐�̏$�I*(Dӟ٩Հ���94����-z�;� s�[�o��>7s�*0�z��s�"l7�:�x� U�I?;���y�L�Ɖ�&�
~�� �S�­D�u*�W�D���[}�z�2砱�>*RB}��7��\��˫�`l'�I��߱���(^Ű}&W��$t|o��G!�5#�^+��P�gb'�ٞy����o�4��`D�[�:�5�׍�3q�(P��ƌ�5�|��\��fX�� �?hpӳ>Mh@3��ƺ���~①���t!4�e�q�tJƅ�݉t��Iyq�.{����ў	�~Xx�fZ-|纛�?�p�s
y����mJ7�]�#�`H�1K�;z�W|Zn�z�t��)���|��
0��S`Z=� g&Gɫ{���H�u]-d|�G��^w+��R?�<��BP0bi�"C,{��Gs�~��sQB ���,���×�=��R�nyᣂ�YQw�Ցa���R�ˈG��h\Ҙ�F�f�Ս�M�ܕ�;�����૖d�c�I� ضQX}��?��
��U6D�N�I9��^[d�"��׷hg�k��:8K�ӽW������BRT~"�� ø��v��-�dta��2��KNW:�����3g� �k���y��`�4��qMw�܊��B�x�D�5t���xX:��x�5��Q0Psy��Ԝq�oZ�~\��8���� ��^���o��=�&��Q1��I3�徎�'��x�����}�B�Ϥ��^����N��@���P�z�86�#��0���o�w�+���;Nؔ�#��,�iI��q� ���c�U3§ ��D��s�,��o�b�j"��1E��{�")b�I����+� ܵs�؉ ��p�2����
��e���>vM'1�7G�5I6e�)�sx�AGW�a (���*i�ZD�do�.C�H=a#1㌸M��N-;�saj�I+Ѝ��6��[�FM<|osR~
b��Z��?��X+�P�c�z�^Ԧ��[�J�>��k��k�߹�b�e<`C�'�����j����YhU�2G� $e,_��~��J⧜�����!�t��?x�C���;ܶ��ϰ������u�`I�o�%��XQ��9v��9�\/�J�pB�d���:��TTY9�U�����.B�Lcs�r��j��`�.�ZS,@3HD�N#F�q3��I�u�6p��2
��WE*x�AF�,�,e���^��n�]2y��N%���S��8���y0(�<b���/����.��8M)��U�E�⾜��r��^�K@f�9E�A��8��`����[w�D y�e�skp+-����V39��=�d��\� c�	���������t
}&�.$��
�L���qR� ����������4� [�Q���jq,���k8G�r���	�ߜ(h49�{o���d4>7ae�%ׁ`�ϴ���1� �߁�Dס�},1��(�O���ik���[����?��k�m]%�7�1ڪ<���U7��&�s�7�4y���2�׹��ҍV-*��y.��ZfZh������ƺ��yo"2��W�H_9W�L��2��Ń�F������u���W��i&^�	��P�&�(^�\�l�.���Ӂ~�G� ��F�x�>pA|�Пb<6��?�rѵ9^.�
h�;��F���dr�?$�1	%Fw�S=d�����x��^0�5�92fs��3}jOK���/�ɑ��0�9֛��T�\)��y�����&�K����E��Ni�^�v���6�_S��G��W��iX�]g�]Q���aA�q�&؃*�#[~Y1@t/�$z5|M���p �1�﨧��mⰸ��	 b�e:(��Z�I(��9�w!������^��ύ�J[��T��}bƌ�PVD���u��
���nm6C�I�S#��Gl�$��Q�ȍ�̜���O�3�w 3i�&ܨ��_%<P�N��aQ��9�::��Gǌ�R�A�Mɮ� D����(Ѧ*-�����s=�a R��_EWu��`c�u�	/��\�z�= ��5�*�i�LsOc�U�u�0�b/1��p���|�t����o[�;�J�u��"����w��_տ���e���Ϲn�@�s��4?�o90;�"r�X&�7��YM-j�T����T �h��O,!�y��q�w���[uT9��m���Q����XzHl�j�%7V�ڹ>Z�4#�s+0���_%���w4�
�w��o�&��AS-H�bJ7�u���{��Tڗ걬K#��O�8+�+��_³p���뒱��rW�L�*�������^�Bj��ݎ�Q�P����Ҧ����w�����1ƍ�]Յ�R���Kj�&�S�ܣO�g��^M��x��sI.���'��P��MDa����I����w�+4��Od���T �B�I�χs�����B��e�5����z�q���1��'Up�i�_�Hl�����o7�;�g��}�>1%!��V�?�	���4��$����\�VҔ��X�:]W`('aӕYd�ŋ	�]�ی�Q��ρ���W�7]LJ�C%C7���˯���8!`�%ڱ�_����]�25�2�˃�jy�]
��gO��Iϖ4$e����C��no��z�nP��K�Myo}u��q�S���ߚi�d�3Zt��R��WUy�L���	��� ~�v]B ��un=�|�<�ʗ�-_���8�B���g�>�C��̀NL�ʬ7�H��wنz�����"�7��Խ�s��"9�X�����@���� ��1˺�x���͵��<U���OX`8ѡ�ںN�ђt��Hu��25��������+�;��yR'Di�}�����(�#_���"@��5�Uz��;8��U���W�.ҔF��.5lƘ3�Ia��K�.���>Yf���B�N�~����]ک{�P��������=2��[a��:?�Bgg7�qZ(h�Uh3�{�%�Y��x��I�a��RccV��z����@y�'+��7�|S�%�h��k���8#�Ŋ�0',h��
��|NҖ��V�����f?Ru{������?͖�|����= ܽ�g�̬NJ�Hk��%�[��A9�<ew��.L�D���A��0��U(�����<��27M@������1����R&��-#�nk)�t��&ꖚ��Ƅ�h���MG�|	u���IQNgB�f)q�C~0f2x&^[��لjMْ���ܸ��v3�!���u����S�0��%Z�Ϗy��;L��+̉�r9�0�~|�����E�J;�
�����(�><&���[ו���p�#��އ�X��q��T���;3�+����:��S��sߌ�Ƞs�m��G�����TA�zE��{n ˪lo�ϊ@�ҹ�ݔCO)A��dLsl0J�v�D��ټFJ���x���YRT������B�2��N�bNP>��s�9��2h#��c
H��cl��J�����֝����uL�/|ƋB�
7#�hQ����Go5e�h͵��/9�O#��a��W�_�`�H�K��=��@X�"
�s"�XJ8Q��(	��l$����hn��>�&��ZO��܊1؜�� �ү
i5����� �ZP,�mu�����dP�3�T�[h�f�+Zl(��#����&�2R�2w��GTɇ�8�M�K�dK��aȵ� �R�IS&,��K���Z��`7	2���xZ)�[r�p�k��D�9��,��\�SO,
�jv�pK�i�!�g�'���4�t��ĉ�,,�K����b��=t,����ä�c�������L����(�~7�}�T��/�������+�f���q���I��:ԛ�ek�8�>`�����@�IQ"��{���N{P���֙6 �e�����%U����S�g��GG���>�N,���e��ZN�k�ΰ}n�@h��}�4?����EW�4�Ed8��Ek2��OVh�1%;$0��[X#��-b��I����sёRs��WT�hn�;ۙ!�:�@����A�q��aen!_,k`*T�i���7�X}L�اMh�AW2�Mvb�¿S��S������Or�L��Ȟ!]�^�<���?ҕ���&���a���v?A�}l䭘Mgc� ,��5-^�*�����>+(L0��T�!�4��+Jr9���B�v�d�%0(����?P���rl�m��E���N�ٺ�*=\�Z��!T��%�����@�{����=�U��RޓA!�dt+l�s�_�d�-��j�N�J 
����LW^`�i�@N�$v�O���|��b@V���n�X�0��I_~������Ca�S�T�
�@x6���itDW�C�5V���6Ψ$8]Y�Peޮ��RKߞהb��Up��k)�3���{���	kN��^���eiG8�����"{�I��M�����t��=z�2%�㊃������d@�ɦh��u�4D��s�[��UzX5В���?��d�C�5s�\�����lX�A�rB��_������j�i�F�{�s�Y~|��
��L��:�|f�+/0Ӏ��B0�l@@����}˪�{Pl�ۨ�E�Ƥ���s1��e� ���_��8�K�v����ɝ�/<�]�F��pU���LͻRUT��!C�f�ah)�N����G ks螽D�<܄�j{�r�}��E1v9SS7��2�ڎS�*�;g���b��.� �f;G7��g����f�������Px�+0OEz�Tj��`�,���0��g��4Bg(�/�l+�[��k�g�W���pX7�4���BCɝ�'V��:�Q{��\Q�<blU^!PaL9����z��A��Qp�k����nNNS{Lqw��m��	���@�U6���'.9~��~4�>+�k����~H]ჾ�Uwg�&8��i��F��AȐz����Xq�r����1��*���j�Pn}�N��7�:I������~eXCD��Y��k����DG%fn��M(F�2�����݈��lo[��Z���P�(���*���Tʹ�7��܊~�� D'�K���,B}��eP�s���	�˟���}Vf��[�E�
錝!��{�g�JT��������НWz�o0��5Ma�3K���t�II��\��T��3Mu%�.ٗ��تr�Ͳ ?><�Z��K�J��|�|��3HG���uN�㊴�\�Z��G�uU�F���c�W�=Y��c+%��#`��p���E�rí��E6)*F��p{�gQ�79��y2g��Z�����	���	�ŷ�J��0��Ԭa�~+摖U6��~D:f�~�<�҆q��]N!�t(:p�L	�}M��m��r�	�C!W��˹"C#^�Wk���T�t�&��_A�:�2f��Z�5�`�-
Gg/��D�D�dykj���$B��d*'��E�Hx�  q%�9�*vC��{��vg�h��Rgl��r�6%+�l~P^5����n���V�4���3+>=�I'�>�̆�q�ҽ���_k�V��y��t�����^3���/?���!p���ޣ>�n>�b4v�j<��zi�겴�T�r�į��P�n��;=��K202=��սs��� ���R�Y)@I?�%H����G���<O,5{v�#��j��{oȄx{��d�]}JxB���Y*���L��\ ��/2�n"^��\O���8向]�5��V��'x�D-�3T�ё��(�ͭ�}Pv:�V.��n���BV�������� �-���ز�7M�G�H]e����,ԨN���W�|�$�G��pȡi��X5LVq[v��|�Q�{���|��8��UG�)����j�xם@Ф�>��$X���.��9�YG/�C܄�J����p[2�l��Ś��,���9��T�t�mA7��u�'�L�q��Gl=L����#��IK¼�Y�/��G5�a%E+\�D+�+�ݏ��v<���<%%�u�-.k�-4����������E�z%a����c�5�ch�\��x���E �>�,��	`{�3�> ���E:'?� =�,H�e#&.�4Ke�Q�8��n�r�$�T��o��v�s�?����a}�!��t��U����M��� [�6kg9:ڄ�Pާ��Ϩ�����+\Q�qd��	U.�A�J��x�Uop5w��ÞG/'X�7�V����6�3g���~�i���ƴ�DG'+Gw1��&�:�bȶ 7�1U�BF���W&���G>��]�{�+����h�����|L �1�ā���FG��x��V��p?��Ǒl|��478*.1���ij?$9[��G�h���Z�W{�#Y��A��(��\d}�(7gh�K��Ƶru��i{O��qئ����cx����ɩ���o��beP=l���4	sN�$�U$#r��)k���xФ���[�x0���d`ٻ4�l�sM��4#���R�D��!�ç.v)��ݭ^BĜ�O��ޚ�f�)B�py�\?�������7E _j,���3Z9�%���z3���i8�#��w:,
9T�0a&����IL{�}�1��Ka��v��»�ܼ�ZR��'�j���z�sa�����i-ɰ�δxf�DȎq��}���b�e5�Ƌ/x|Z���cF��,�I���gk2���!��ڽ�7 �`��9a��LS�BZ>����2��·���{0�=�r�kl�|QI�!e�zы�
D�/����o2{ެ��)m9�:�1��^��!�*G��3$ô�s6A����eս}[�����U���M��x,z��]T���a�KNb��9 xB�G�����=ȩ
���E�W*&>����<�G���FgX�K��grc���$~#;�R��~eǹ��p��6;5�|�vc��Z7���$����4������2]U���ï��	ً���p��s��6c�ȕ6��ϻ�(a,��F���>���@�!>�,p�W�Z���b!����m��3�A}vA|F6��������+�T�܅J"T���ߞ��EE[����գe���|�#�B
�6���tY9���)���]�������z����"�Y�!�A}�SA��3|�E��L+�����EU:�s�À�4��7��=܁��o$9+2{i"�<�|���[��i0�ȇ�9��͢>�%<�M�SO�^Lv�hF�yQ�R��A�#&?����D3��
V%��P~2���<���N�8^��Q
#D�D�!ZX1l�������u����`�q7�T
��T��>���]�L��d�Nbȴ_ �I�!s�W����#^_�`�zl��Z����e�R�$4��L%�dx� R��h�;)��ڳ�#hC�Dd����1��<A�Y�P*���l>ZL�,���r��S'^Z���L��,�6�x�81&��+a'<��*� .��sX,�P��m7�)����>+�I�J
�-=�6�!h6����i<��/�M�L�n�Z=��VI�(M�2���mA�oM�&t'w�^�$X��iy�)��$�@�<�#�(0H��b&8�9Z|�&왜+<�E�f.a5��2J�ny1(���`��������ި`q����t���+[�Xw!Ď��z�y� �3����Q����o�8}����?�OΙ�S�qѓ�#t����uWѦ��nq;���&�� v���羾oP������*<�x\3�}���3�3>�5i�m�
��O�S�f/a�p5`f�+,����ƞ�Ոғ�A`p%����%B?��&�>R���qd׻;�S�321���Ǩ,�{��Ѿ��:�P��u�?��Ή���(���$b�f�AƸ��h�b=[�|��mW��w�v����Y>� ���j�6ֹ���z�s�c�H���)�'8�hE8;��G5f��C���B�#c��F~id������. �|���vp-�=�]�L��ބL�����g����j/��W�8;�a�G����y�7����$P%�^���	���57$*o��UW��.bs\Zdl=S��Ŵ�ȴ���2{�)��1S{�?xX��� ��V���G>�ἰL�f�z�!s3���k �Td�~O{%�è)�1]L�q���I��2�v,E�~��-Zެ���s6<3�l�~����l��K�"�r�,W��nx�jw�Ol�tw����j7[F������I�ؐi����]��+���U�����.\*'����L�Ke�}�c�(|�uUI�q������Q�y�˙�Z��$�OoŊ��r���0 I�hm�lk�@���;'����e.�iKT�)��G�=%W:_W���~NU�� �I�5/�e9��"$}D�{��9zZV�Y�V@������u�C#�Y<�����0x$��O�񇼬����<�T~�~��gd�!"u�U���� ջ �	Q B�������	v��ո���}S��{ؗQN��J�m>�U?��t���)�s�9��y���=RTwm�w��n���$�5��_d0D)؋h|� $v��)`�h"R�7$�2M{U]��h���E|]f�:_m����]*��Sg�S����x��>Nvp�{�9mD#NV{mp,!{F�jP^dH���l����-m�@t9�f�N��E�zRW�����c�ƈ��P1�^AǿB���ND��d=�Y�~�/�Zω�X/�<l��!
�F����s�w�������!������-�b�$Р�y�pP_� �Rh�%����D�O����xaE� �a�ɼZ!�~%�R��[�F�ҷXDm��|�a7U�]���sSi�p#��K��]^Oh9��-��F�����]�ι��� �=�"�>X6�e٩�7!�#.Qe���/�� �$N�WI�:��ӟ���xc�� s�>�v���W>���ф��& $B�$tch�*��&i[�}E32N���yS�lr\�����nK&|�%N^6�^D�2.nX��}ZD�C�<����4ʞ�S6X�������;Z�_�9���v$��O���a�M�A�"����	M�D��+V�e��W����)�7�2+GJp~�'�D�幻��@�r�4�ƃ�pR��$�Go^����v#w��d��Y[�g�n\�;��$�?jV��� '/�p�.1�p�yUa�x�Ur)��oD�;K��y�fTN�ń��H�c�@�4�0	X%���XyCH��CRȖ
�E	��*��~���gرaU�	��5��G^�'cB�?�����(�&X��1� ��i��I=6���c���Μk��dS�Z���T7�������
'	d�-����X�ͧ�X�4<F�>�;�x���l�p�l}9�������Y�?��IX�HL�Z�|�܋O$h=3��}�z+��#/����իN�ٴ��I�PDQ@�.�x�՘�m�
�J����-�܄^�%�����,�L$�Ya����"R���Z��� �|�s3��G:<[��[ڵ��0�\4���W,_F���Q�vWB���X���7p��.da*I�y�������5h,�˨��D�j�s�3���8�d��uK0��h �ro1Ĩ6�����C7��u�}Z�d�F2*8�fY�2��Un�	!A���X��~��v�����>���o"��*ז9TyM|J�2�H9�9�����KՓ���Y\��
����In�"l�)y�9��;?a��z͔kh�~^�V��lt�����^�{��,��6*MS'$�#`URAR�+�Gr3=��K(�b?i;���?yj�fIӑp�xiX#�z�������� �E��|�j���Ա�r��=a_�b���X��݀XUK��O�{��v��ዟ��}�:���4Mc��Y� NV�J�!#�07��zB��I$�0Q�+$�)�P���a��C��O��ȃ��P�#��]����������n5wH�R"f��,��~��K<FL�_��H�Oc�~r�ـd]/�u@2)m�8��k7dkz�_�@xDKR��0��e���j�+m�{<F;*!���LB9�R���B�q�A���r���	M����Zң�x�V.P!�>��jq�\H
�I�m\B��Be�x�A��Ә�ڇ�){ �^�U�d�X��,��2@Fi�"7���(��5|�C�TRѬ��6]	Pb�J�{��0 ���"vJ�O�4
�{I�GK�/z�8|��	��zE;j�$�]�(��U�1	�'M�M�Rr�k�����xgU��874��~U�5�Z�_iE�z��Y[p(��zx��n@��}��i��=���<�i}��2�c�����[���r�)�Q+��*U/P��������ɔ�����T�R���4Y���>@��)_1��^�y,�g`� � ��=��B%5�Mi5�C ���J�0˰a0{M��|��OZ2F���k�D�]�d�K(H���5���\��.	��%�č��(�D��=og$�[*�+�-40V�$�. ��T}r�өuKI�Z�1٤�p�LƋ�8��U�m�S�:�,1/�.0}�M��S�4�Ϫ� �����f �BF`d�F�t(�8̊�vsȟ4��8�Tp���.�'q��8������dD�f RO֢�?~��U�?_��`X\5=ԼK_�dJ���Tk)oe�|u԰Cd�R"�����[���D��b�)�tD�| UZ������2ٳ)�:R\�"�لd8#w$0��W�߫��F&�� �f��΋����Y�@f���BƐ��C���Q&�CF�7�nY�!���s�������D<���ӆ:�lڪ�5PrAoŰyX:��^@W�|@^�k����Ix��.D��	� ����j��PahG�Y���~��/g�,�Þ��A��g!.��ژ�c�P@f�����p�h˩	a��M����t��u}�{xc~�C�iQ����벏�L|�%��̍C���z�<Rǜ�\�	���>U�G��^�Z��n���\�$�c����\ĭ�/Z�<�|B�Y���,O '7�`,����ζ+�"x�K��a.���Z��DM�v�;L�*�g/t���<B4Oj�{��y-��݊��Uϫ�sd՟2�'�c�`*>�,��x�=�(r��u��{��.�P��nTc�x�,0����$�\y�"U��"q�S��'�Z��бĔP�K��5r��	~+ed\����H҉����/����Om�'�u�q1a#xc���~���
թh�Vt���g��?��xv�gie]Z��9}�5��:����{�~�Ef�����ZfM���e�1�v��Nӟ�{�ݯA�i��
���$6"�@��z����T��Ȉ����7(ۢR z״���l+G�?Ԯ�<�9"�H�=�6Ӗ��?-u�~�/n��o�n�5����%��Y��?�v[%�' �e�'�̔�u�.���)�b�T���D�\_��{��"�t@���"�E���=�϶��{)���6�s4��q��|e�7�F���&ֹ�U�� ��t���N�ɒ5 �'�
M�#o2�v�����w�Mp۾j`�g"8�y�$y���>wC�@
ʺEo��Y��#2���\h]�h���N�6�}��Ub�b����A�_�gW��{�8�Wl��X))c�H[�W��L�A������Y�/#>�0t�������|�_\�	���I�-��q��&/��I�d�O�+f[��XHRh��2D��h�5=~9��a��"���lu�	����Y
c�%�xQp�d>H�v���X#���I��'Z/�6�Y%���ǧ�P L͍�_�j�/����Al*�]�j�u�M���1j�Eo#GB�X)���� 3��g����5�KS����J�(���5��$֕�7`5��	�~�g�����������I��q5��ڵ��p�����/{{��&������mb-��f9t��f��Uœ�$�p������Dm�����F҆\��3�\x'�ŷ�k%�{�}x��_AGO'���f�'|c� �PaqVSf�PY�H��8��7��YZ^Q慑dfX����^��e�������,\�j��sJ�������w�r���Y�غ�;P�<��s�,l�⪧0ЛL�nm���>Tb��C1�R��$]x,X�p��g9�JJh�1�̏I�b��	7�$�ѩ��q�j��W�xbA��"c��lĳpѦ��E3C��y����`%��o�m�Ϙ�C�qdދ�ma۲��C���e~y�iNw�U)���\@���H�	���Y�]�a������t��l�R`$��j����G�NA�՜=�a���,����������i)�_K7��}K˽S=�.�,�A�����:�GI�c�__�����SR�oa��;˒������l*Ϊ8q�\����S�&O\cw�u�!<�� �V8�����Y��?>�@D������]��]4�wʦQ\�4��j4�@U1�~Y�������W�����5�ε��T���B��w��Yo��?8�m]�@�
⡺������:�m^���&o�	\��Ǒ��i�?=��Y~���T[LF�`�3c��t��"�Ne4�Wa'*��hXG�)����8țm:œ��`���e_��#�J��*���E^Χ�*$��	��Zt^��F���������W�^�SK�j"��X�<iH�*� @� �����Kk^\��Z�4O&ƈi�v7u�}$@���&�ɀ��1�m�qҬ9���Lr��d��FpuӤ�]���8<q���U>����{ۭoV�6�`[=��ߛ����Hf�s��Yh�>�	._j�iuR������{#@$����R]=��y����>Q� �Ф�8�<��]Nz?�ڬ��gT=���uW-��5�UYu�#{8~�+a�d����񷎐7Ȇ7�pG�|PӼ�e;y�zj�FM�FP'qJ�WC�*�y�$Vn!����Q���^����.{Y^��i0���*���2Vďm�_5�x5:��B.�餇c������^R�r� ���=�eCE�Nf�Π_��?N���6���W�*��d7���D���� �G���v�DA�B{��۹�J�ٕ/��a\��ɴ��m�:���ϷۏI:�U�����W/��S��R���j��ʛ�O3�NǼV Sm��bݧ���\��o������H�R��_��E��e!(�R��'#���ae�1�ωcr�5�5�<���y��i�����j@
��͸=���[��^����u��������&���s�7�J�9q�TiI��_G )�Ję�zަg���[��q�ԑD!��U��C�9�:�4�^�� ��ڑ�'��ĩ
<P��} ��A�4E���x��y���4���Q�V�����
�v�i���1Թ4��8����ѩ_�a_+p򶂦�}�-N�P�1o���~z���rE�<}e�"=�~�tV�x��	�N���sf-�^�����O��G{?#g�(B��D)4X �;~��]�b&��$�ߋ��Gͅ7c:�.�ʉ�N����U��K��v�<���|'z�{wBCX5����-\>�r�}c��K���f����7\̒�Ұ�Z��R��g�,Ӧ��ȋ�З���N��k`G@�U�l��7�f��;Mک�e�=!��r{��.u1;L<~`J�W�d�CeCP��������oz�pу:���>�㤶ۑ1�"��ë��l�# �6J�wq���ѵ���%�P�L�e������@䏿Qz�[+��ê��b�mW��6�<�:7��\T�u�2R'4鈍��y��ϖ0t�F �SO����'����I�� �E-vK�t�{���gOiN/�ɕ�W_�z/� txJH��!=����� Q���:�:�Sѡ�<����G���3�o�����Rq}�b�f��!ڏ�M9� %��S���Q"��ғ1�竁k�(p�J�2��v%�����}
���(s� ��E��gr���,����.D@#�L�>�ޚ�7'�/�w����_[H���2��x
�bM�Ҹ3��n��[�)M	߬�k2E�����N�&n|��$) z�ȄA�MO����[>$�=�>|Q���K������h���k}�DG�]Ƨ�<���~��'��cy����J�x�ގ^�����	�S9^և��Bh����%F%ߊ�JF
�A6r8���{g]LU��fu|��d=6�$�ػy'8A�	n7�񚕥�d�#���3�x��n�@����}7�čiE��	���u/�~%�-�F �����!��5:�6f}�G]����	��G���2�˭]�yVzm?T�IZ���91�N�{-�#�((₶#��S�?���{�P$�\�D)=��-l�z��ժv3L2i��;�f���{ �J���N�)P[�*&�k*s����a�C��T��<�c}���ӂ}��5�A"�
*>��X*��َBl��7���N:Ў�8P�f���9���憎�yZ�D�Z����J�cs�3�Eb��M�+��f�{�WR)BRN�.?Dp�`a���h�f���R�����;-[0����#�Ƒ��VWMl_���扎���Y�I������1O%�`��2�R_�-y̦�6<��q�E�v�F舲�u�� ����]!��FF��=��1�1���w����A��#Y�\�����^m�'9�)5�|�̥�\b2�rf���h&P�q�@��v٪t�q�֥�1g[�������ᓪ�.@潤����E�Nd�������rRr�bE���%J��r�b/��W�ڮ�� ��m(��0bj�A�䆉�S��c	�l�=���F�I2
��{��>^�04L�eR@4�'i#R�sVMe�!��� �z���o�L/��f cr���Yg����G���%R|a�<9BS5K�����ub�~ q��Zw�m��զH�Ю-�#����)�C��\����R��^�Eq`�I��=��ɖ�i6��ҳ8��U]��>��-��=�r��-�p���b�L~��7�N<�U�D �u	u�4���w�����
��^�i]Y����PUrR���r&_�kr�,�K+�,њ�������{N�sz$��2ҩb9cW�ҝ�BUl ����[��AY�0��4����'�8|�!f�^6H�����0|#>1Ycĉ��P��*-3�_��;��3���'��T}xԥX�%�b�塑Qy�͕�6�j����ݵ�j��kf���qo�%�5H���p�<��b	Ec�z/�ػ4�^�xۗ��TbBS����y���S7�R��þF�Q���ܗ]<�-���tY��E��3.<�B��v�a6Yd~jQPFe�Ψ�Z�V�՚<�ͥ<�L����24�H<��M�����(9��~	�!&�S�4��.�A���"�+��o��|k�@;���a�WP�! ��{TQ�k������:�L�Aj5$��7�����|��w������[�g�'�U��f�gO��@u�j6khz��a�Yv��_���KkX�#æ�[#��3+�"oe%��#�.1����ǁ:d.|S���W����R7�D��>�F%n�ho"�\��d�T$>��r�%(%x��c�7�,���p�:�%��z�,�n�-x��Z�F���iu]�}��	�?�,.�K;`���ߪH�T�$�X̏��#�1][��ٌ�u�E��b'a�
���D8.��������KC��C�;K��r�����M���~�Ƞ�olPS��٨R��X*h���λ�&u6
��� �{y�����1���.#2���5͑P�1b�>cq�b����Vu�ws�sk�{[c�/W���Ұ�����,�ZL����T����]2L��7�ӻs��|U�^)��l�aJH�v�q�G�E��Cfs�u`��1KO�&��nݬޡ��y6^ӽ�qA$a�	Z[��:c�S�C��t�]^$������@���qb&\t��SBD�yX�.�#5`G��9�D�25Y]�u��A�X-2Ɓv�2�re5�~��beFۀh�a�S�H8����[�=��� P�y��O���]�� i��/p/�v�����2=���_��s �*�c�vF��0� �����^ՙ�B�TS�ӥsO���m�R�w-==K�Sn�7��go�dVƳ�\ݰ�ʚ�4� ?"���bs&��o�ܙ3�ADd��-����H+ƀƆn`������|/�Y�4v�*�����pҢ��CZ����e��*�%���>��%B�@Us���}E�Z|˞	W�/�b��=��5y�/Τΐ�]�NĞJ�y��5ي�f&���j-��]d|y �k��*v����&=��0�bƬ��%��?����E	�
���d�����_���g������u����2Os����F;<y03�|���-%�fg�� 8��!O���X��fj��5w�u�3��y��U}/����|:0o,*��^��.2�>�^�ҧ��5:̻Ї��`'�>2^BP�?:�R�I��=�S�x4u�z�%2��V�������V�_��Eo��.��;5]oe�cIq��cڅ���z���V���w2ڙ�s�T�'鱵/�:�+l�)oH��?��M"�]�j�6cEc��>ѼG{;�1"�9N~�I8��;`%9��3�-��7�bc������|�@T:M�ʵ�.�Si$w�+�������\�g~���=��g��9�k��\V.��%�,���y�f��`?��c����8�C�����̍I���r�R���\{�_R�T��<�j ̏-��\ �:��걎
��#4(��⿔�� &���У�� ̒~.������|�=zح���[�^��Aѣ!Xd�|9�Xc��� �C�:�rZ!
�R�]�w���G�L'�b���ҫ��]������0�gPb����C{MYd��c�^�̳�ܰv%U����Z}�oK<����-��λ㎡F
+UNЂ�m
�����\�@��*ݟ�M\�9(��/?�v#S�~�����Ni��2� M�R���QK'���}���r(�G>*p �����L� �`%��Õ[���nE��y~��j/5O|A�7�����9DT(rm���0;���^.���a;���U��Ra�%�˹�/V8c�@y�pV��V��f��b�'�c��P��n��.3ޔ����`e�G�W��p<�h��@�s������	��j��O��B]�ا�<�z���`������7X�Zm��ꅇk2m	�"�bmr�rV��܍)���Z�;��ArqB�Z�A��7�SV�&S��C�ێ&��2]��KG��C� ����'�y����W�=��M-�e�
ޑ���@�w�D�������)�dmѷ^VK;�^�Y��ǦW=��W՚����a;��;`vm�9�w����I*�zކo&������t)�s� �K�t]y�n3�������g<z���������S���C�t��>���w�UBW�k���/U�`)v8�:}��ǐ�-�\�����{y?�M��6���`*0�=]-�A��!��V�_�����!�i��>W�JΌq� ��jM0[�L��|�r�b�^/��N`[A`��s"�e���G!��#@�-�XZ�7-��^i��~���VA�L��qD�)9�>E�;|����_;��)k��H7�>��C�.S�SG�Rk���޴@_,n:@a�8K�<�������&���?R�fpF`��v��N�4�oQ�������2�iD�gPN&}�Q�+��$��}�+��m,>@� �߷��?c,:�C�\ş�˶p��M�/{��� ��2 �9��:S"��t�B]e�'���vr��X���VH���y؍��l�855闉�Y��&:�1Hhw)g%ܑ��ؓ��2J�2R~+u���7�T:��"9�N��N�e���o�3��#9N���; l�&+2��?����b��Y�3������ug+z8�{�:��m]]h�r�'�s��ـ��GR�S�����%�2V�(N���"ƘX;X��.������kN R�lqK}�d*A裙��"��?4�t
��y�9pzJ��� @�`A��@�χ
̯�G�%hS�J����YI�	�\��� ^�h�~MuIm�A���6x�.���+[U�!�ڃ@v����XԾQ�tv `j�c���j�jB$1

�_!�%m��̡x	ZT�L�tBig��2���.�i��"|Ux��Gx�ܒ�YU�ua�)��шg��W��"��Ǚ�� Ȣ�zv]����5!^b,3A��J��lfj��B'�����ku�Ѭ�+=n7*�G�Rb.
�'9���G�_���%�BG���4�6� �H�{�4�Đ�!���WȥҜ;��:�&w����aߵ�N���`�%�����?��B��MB�8(�,�$��dc��򌥄cH��'�x�����F9��$y���"ֿ/���o�W>p��N�)!?ʌ �j���S4c6fNg��?�V�������ig�n�j���>���lRG!זj6���H0m�5�n���@��F�V1I�<<O�6hֈ9<4��n�u�������/�t��V's��Dd��f�؋` %��P���V4�*��
|Eeg�$já�%���Ӂ9��f���ٖ�1�NJ㏼%�b�Ģ�)N������/��᷆�ѓ}B�%kT���o�����b��_$Rwq4V2��rt�A���^x�����(C��{��<,���d��pܕ_;��$��@��7򎢦ûB�a+��N�*|�#^��O.�=AA�p�(:�E��UuSݴ��b脔ʬ�+XǚJ��D�` �V�R��!-�b�]�qT2/���]l�L�frߵ�8����
�n�zU�G��v�0�l���b������{#�_���
Vö�E��|:��$ƻ��DP���XlV�/���=���`�	|�9�_!��٦]&.����h���vT��Z�Z�LAGAE.�������7��{�lqk��q���=��WǦ�,7N��Q���5>�<\.qk�sR���v{�A���Y�R˦1��lUy��o�3�V�|#̭9-:���mX{�oK��mV��d%>{�����pD�P�Z܄�3��0u'�Zd�;�%���Ro�kr��]�̹Xo���\;0���P`�WJS�}-��$�x5N-����i�@�R�1S�)��]:�����BJ*�O���Pr_�o_ŋǑ�Ph�ҳ��N�oH�hm�����H��'�����Ж�d�B ~Y���I2�U#�# `jRC�GI�P����1�o'���1��L��N���-6��1VB#W��G2ilds��>WΕF%e���� �K��+��}�
�jP�u!��Y�l$5�Ȓ1=����ڜ2�	t� �z�?Ȝ{Ҫ`Q�C~�w�^�6�nvq	�éI�wݠ@[G��o�+��d��}��,��^�lP0[/`qX��s3�{�6��m^�	H�eV�`�f��gE��aG<��2y�������($\l���ȩ�~�"01��b�b�Q��h�w�wz:��-F"S����^����2�~��J+�����q�R��g�_�}��g��6K�P�w; vtR1��#8�2��#�oC�/�T�f���ZEݴ���w���cҵ6;�L�Yк(e���zM�ad��7�V�"u�J�+/�C����i<�E�r-��va�o]b�[�Z��ɏD|Q�?z/afר�̿z�5�l2!���}?��՚�2g
��Ol��fL��?f�8��9�;���zrG>�v�����P�?�i2�_!���|� �U�D�u��-R{ڬI)�[��LF�b�?M�Vs��Y�T� ��ϔi���8����#���ND�����,(�n3C��^@���m�:�o�$��ۯ}����rk�Ci7���5���Ѓ1�!��V�ˤd�u�{`w�d{OQ���v����֙����X?@|v�w+���+?���8= X|a�GO�3=�7��-��'S���� #7n��3���)1|��\��A�"��J{�����kNWQg��!����e��2����/�����0FR/ ��E�t���� ��=
~�,Ȁ��]��ֶ���j(ށ�9�^(D{��F�f;���(c}ǒ�`�&�}�����t6�h� wj$a�xuP(�x�4#���B����|���_D����v'�MEڶ�_]u�T���&�b�D��/��ig�w[��h�	S��`N�ZD�ۆ�9 9'˃HD�a�%��s�Ij��^�����n�!q�* W�;b֗Oa-o�栂#U^r��@�9����Wx[��%���V�?��yB��q.^'wVPDw�+��U��֮=w���;!�JZ��/&��&�:7�t�9�x0���١d
�t,1��r���5���P6�ap��?���{&YP#U��5��A�ԗ;+��pa�� n��I"�����"��1�_��L;O�/���������#``���%-���?�,,�lB�\�h�0�?���{��	/�A�uUbyEFA�J8�Jͷ[��;ژY�l����҂Q�5��_1G�"-��-���҉��>8��;������~i�*t�x��������m�r�(�����)�O6����Q��g�ew���
(��Ε?�@X�Wokd+�w�G�5���*���!��X��!}��bw�ӭ֎1�7"�Ƅ
��Һ�m,��7`g*"��&$z��!&z�CI7�i� �P���0��_��2!B����l}C�9r�쇗_ñNK���J�]+h��)G�Tr� G��Eۚ�����|G����Ś��[~�}Z��^�(�N�3=�� �2�s��]�ЛR|4$2��n���M���xkC���kѧY\C�MH
E�+��t�(%�f��o����5Du��3���J��3H�s!9�}T1����oe����}�Ò��v4�[�u�gÉ�W�N|DwO\kZ�d���RNf��<%V�	��[�Qc4���k��X[Fn�T�=~
�a�����WB�Z�Ǩz㺢ŷ����)om��TP����'鎎�U'��`gF��l��CX��#�ݮ�P��B�
T�Nf;��&L��ǿ/�1W�Abh���z�|>���R�F.W;�Ҭv�xz��t�g�O��^\�7�jhv���d���Y/��nKm]�ڒ�����7�l������ixnb\�y%_�\@�K�7/]�{���?�sN��9{�
 _F�3��3x����]r�;�z�
����8�^�\&w�K�ְ^�:%�麔�mP��8��c��^�!����p��VJs���h����9��9��;ˡ�V�g#�n_�wT5Tc0�"a���h?zgFG�g�{����Jl�pu8�W=��S�#=Y�h?3R������0�����IJr�b]Z ݩ�t����}��ǙYR����N%P�9�[�kez����#��ܬ����Zk"#�u�.���v��U
���|l$��p�m�@��<fO�sM���ݺ�ڷf�i��~�i�������g��1 hlP&nK��]��C�{\_�P?���PjC]sd��ˮ#z����d�D:*�܈�ef}"�ŔwK\*d\�iyx�)M�?E G��aO=~)@�=Pm2�S��n�/K�G�6���@�q�\=�S����΄�e=(�	��)��w_�
�Ѻi�ދ��5����Chm�l�^n*��w�.��8� �y;���F0q���QuQ�]������~Ag��+:��P�0tFK�4�4���Tf�*�,����b�k|Q�&B���������xn��A����$�R9#�����as��a�vX����.��s���w5�\���*����m�D/��]�d޼{������w4��d��P[��D?VV�U���B\����Ȫ��_��^�$2l�5MƮ2�͔��YR���p��Rl|�$���{�V�n�K�F��J�$���ǯ*�tB�IjJdNH����XS���C4WX�=z�YX��}�#���V*���<W�6`���#��y�;Bb�
��A+?����՛������N���Vb��͡R��a��sP1��W7T&k�+Ցxg��O9��ӄ�qu"^�[���M�.��X-�d�Q�%�5�n���!��h~ܡښ9���n�}�'dbF3@Mct����#��a�1/&b6�X���[`+��p}��S�{��l��[�UK>�_ĸ�ؾ�XS�g{�C���q����j�T��e��k�A}�cM-rmڽ�Lt9~����A�g�0��5B�oV^S��n������CY�#/V�ϨR��JRT����:6��Rʄ�2�%p�=�tB�G��D��.��Re�#<+�i�f�Ӈc����o�y"o@(��c��I�����!����vH2�*�݂��qb��H�:	�T�B�To�
;������%̾�|�o#J�U0(����H:�gӺB��}�$۲�
���9�������gY��j�s�D!��u�!rk�t��z��P��E{�4P�xSڔ�j*������,�o�+m"�$�۟��T��_��t3]�lGN�����ȼ��6��� �{e%�8�����;7|"��ߝMPBI�Qp��F��1���0�� �Ή�پ�Ǆ����BJ��]�Y�/kg�m���,rK�5dagg_:SkN�']WW����g�$
����zNy��I��-8Ǿ ��I(e�$#�u��7m>�P����gu�hQ��5����GS�V��0$:8y־Φ���˧�����t?�'&����;�Y������?R@�S.6 �$h�D�J��&e�zXs.'�,o�=�K`m�$La��A����WeX��4��2�A��2:߁3��(�X�Hf�l�y*)�Ma�	��z��Z�/�����f-`3�{���ʤ�A���K3ү����^�u�4�#�\g,j�_β�5�*ʜB>�
���A{'c��\�Bm��s����h��"g59e� ��/��T��>��cf������J���TV���Zp�&����Ye��"܍:N�l�����l��9��M��<�a��wygV�A�=sf�[����*���qg6���ZLX.{hPQS5ƀ���o�H^��+���pV�ͭ�xШ3>`Bk�hp��K;��	Z�lHD8s�[C�AX��Ayq3�!fs�1d�IP���O�a�Q�:��b:�����)f]�0��ر��Et�20��t_�q	F}���lӡ�*c� �����(�D%�|kp8P�[� ���'��[��h#�����:��T0�8Ì��Ey��mٝ����_�V,D��x�����<d���~���Uj�3����p�^=���n���A2�V��d�L�����V�a��v�&���X�(����r�)�o��pO_N�	��X֗��2��Ъp��i(�~��ؑ��p���a��#=X F)����,g:!�����V�.9��],�O�����b/ֺ�}K$)�5B,cs���c�	R[V���	�3ۥ�'+ҍ�ZVN-V7Ԑ=s�y�P��e~�R���2k��;��9�Sò~��|��bI׳d�_��pߏ�K`�k29��R����c�1��mX]�3"p�����ZV��jz!�־�S"2��])���HHâ���n-Ǜ����t��a�|�2ԛ[�@�1��&]f:Q��O�,X�t�ֵ��Ĺ��	��V�ci?�JO�!s*�}i��+'1�'�7�C-�9(ȹ�(�S�lԄ����4��VX�� "oX��{#��H�o�=���EC|2~M�*��+`�y�D��帆�I4�]����O�n�A�fe��KCq��".����UZ�T���}�����jZ�q"��4v��p��$����ŀ����)L���X�G�.�g��x��ӣ��3�^T��<P��]]�f�[�37H�!��=0�U.Rd5V�*� ���2�nS5���s����=�5k��ӚXL.�x��J�,漺�B���g2�����5y��#�/K�C�ժRҾ<��Z�j�lU���BQh?��,e�7��Gᗖ2��}	P�~�i}0�S/4�W�@�)�O���O�KZ�o{|�ߧ��|Y$��Gبy�Ǐ�n��?�Y&��c�:��&#��*��`�D7a�6p�=B��I��hq�Pc��7Tp2v�%��O�Yس�h�ed��ѧ��H�Y�����Yw>�0X���@��++9��~*9�7�`v>�.J�h����΍9���[� ~�^�3Zt�v��V�$�Ol�n9|��QLMX���g�K�E]	̹J���D��5�� [�Ã��N��20_I�L��>H������9΍�W�D�����J1L�ө<|�U������5Ql~sr� �h'��o���,��z�x����d�|��GF�){@��]�L��.�7L�?�kn�Jg�bW&�u��;p����=�;��i;_��4aگ����6m���{c���	W��o!;s
�� �nb6�Ϟ�jw)J�<�gHa�u�5z�J2;��!�IT!���m�Al��I�pʐL���\�f�f~�,.j#��h{i���]<+�O�Q�V^�1�������T�'#��D��a�Ϧ��Q*h�f������g�m|��	Ah<vN6)l����l�A�7m��@����#Z��3?w�~��D��=�s���I]�ऀ�	>NA�a衣Ʌ~�c�*y��6nQ�~��B0(,���1^ߜ�.%}���C�{y�׿����aMT��R���Y�wYUu�S_%U`�r��!��CE3^"	ί�4;}���*��$|�����_Unt�	�׋�צ2�I���ًJ�9H=���4�hp���d�.B��Ș��6����FR���@#o��È���[�����b'HE������[=E�q�=Kܼ�P�]r�*�6����5�0�j����(E��[&��b�-7O��L���I����ι<7;&�p[l£>}�e#\�(�O�ډaZ^���E���>�(�����X�s�u0�?&kW��9�"��kQ��p�z�_J�����d����8�>���e�;EU�=���Z�@C��������^N�i@�HfD]+g�Sh�.�/�W���m��ʮRƂ��1�8E��9�q!�S��s;C�@5\�F�݄Nb_c%�,���Y"��ٌ�#�<Gk�$P���Qh�N����~�I�&��E��X|{������|�w�ܘ��&��""KJ�ޯ�����Uz���:ѷc����e�d|�0y8��|�u���"�>��`�|�=KM�:g���w`8l���P�c(.\8U�̦�DT��$��٫J*��SB��;%�Ex�K,;a�]�왻����f�����_���wqL�6�IY,ֱ�ֆ�5����{C4jd��=�6�h���`��$�E͜4�#�h(�Xi�:�*"1שO�U��+
�����%�Q�:�j���|�����p��Yس8ө���1z�hy� ��N��)'H�x��b�P�(�qnX^�2�
p�x㋡�oxQ(�Qi���Hn��ԼU?G�������V��G3�~�N�,��J 2$$ʛ�b��l��U�<s�����|2����{������a�����i�{�q��V�a��L���.�_�.C��]K'݈
0�d�(�Ԭh�?.���w͠�-F�g�5�n����;���h@�wy�!��k0�X(�fO�%��.���s�%�$�2R͑���A9-m2t&_b��2�r,A#I�N+������%��I�B�(w%��fq�1;��{����rO}S�$�T�_�Hb8XZI{�#N9�l��T	h�2ʦ������(a��C�k>D|N��­Ю��p��mM=>���M��m,L��y�ֱl�r@d��jڱ�d��7g�*���J���"��L��t�C_�����i��*J3�5螖W�䛼lJN	�P(02���ԛ�lb�=���˃^Y������FL���g�y����Y�M��	a }f��ȘLh>�v%Fg���M��,��~��v��i>Q���юY�v^����nL���� ��1�؛~�h46TN4Mv%_�J�k��la-��H��҅,1x&���cv3�N����c���gw�N��|(h뵖�I�ɿB9<�=Q�x;��Yn<n�_^,#x)�£��9�<�ë/�NVj�ߢG�x��;�����~��Ede��&D��RU�� t�@�ga��JJ���,6��=��ҏ�L�{���-�A;�Ն�{��&��*��H��=|�lnǤ�ʣ[Ub�0��E�D_��s;a�2 ��c:	�d�~�([��mȈ��/�'��bOH�/9�k�1$���,g�
6�
s�-puY9�B,{;w7�?X7��{\f�qM�M�f��N����&���ߵ�c5�o�$e������l�O	��(�!�����T��%�n>/Wu��Z��z6�QO=Ey{�@*W.��y(������NT�Ж1��m؇����A�����z�S)���O�K�ZY�F*2�����%��+_H��N��z��/��o�ԅ>y�s7������y;��y;8��I����F9�t��4�`�cx�b�c�;)c�������jٚo��	�1A�t��6'�7��zm���&��������mD�9�k���)����c2**P��[����U��&���Dr}	�e���Oh��zo_����t����Q����u�_�Đ�Đo9kc�?�Z�r�����_��Gr�սz͊�zT�.��K���?'�.�H�ܢ��,�P�/ء8�W�c�P�9���0�Ω�=o(;���W<A~՛3��2D'm:#�:Ҩ�;�=����THi[�$��`����R�YdԯGZ���Rc������\vU����K��pj-.�g�F��0�e͝5fS�1� ���Q��!W��*����U�'L!�
�镈3-�������	�Zk�s��|���9g�*rv��w:FF��!��7�L;c��m��*I'�Q�ZD����zZ����ȣ�2���?mퟐwO����J�����eo<ю���p7A��䍕��钎���<䳼O��[<&c�L���E���kZ���
A�&,�ي7k�9=R~��`�ui�ؖ�/�W!�ˑ���KW��ZQ��~� ����U*�H�A;X>�3
5LIp��i����Fw'?m�N��H���<�j/����q�;2��1�PĵY4�"[�'���%�}��E�]Z~�P�E�n1�4��W/;K�����黧QW���>VHFln����4/?�{}R`A ���n�Y"��T��ƀRg��ȯW�|\ߘ�ӻ�hl�&��'m��У�v�}����e䥇d�@'8�B{��ۚǄ���@^��@]o�I`�<�'��:���b��'|��cc�c�y�W#�s,�V"��Ϻ��$�G|d
��̗���6L��	A��5�;�T����x��o7�(���Fm���ZKACd¨�&�6?7t�����_&A�]#%��?VJ���눶�wI�dv/Px�������C�.smIp���/M�(�h��(
p�s�%�f\�K3�-��g��q��*�]*_��,<S��0�.W�����Q��(>��M8]�#>U�vN��d��V�y�p�,���G��D��|V	�;��Q��8��,�d���khk�OK��!<��H�1Q!b�����9�wI�b0���!��K����G�$l�;�6C��U�l�(ߢ�z�Hn.��T�9İ�����ou���,��y�L��y`���1)9���M�B�C�o��ۓ�	 " $��	��8�s��11L\P��G���$Ha#N����z��q]K���5<���֎]��FN{?z"���2��y��k>s�^�k�G��F8�����'�D����V�$����!���b��J!�鈕�/�j��a%T��ׇؕ�	��v�5p!+�g!Ó��/N�F����nt(Q�d���`4s�j�+IYvz���D5���.WLb�i�@�H�OI�����x��=z:�<��?(0AVn���M)b����yK��[f	�r��L@�#�m���ƛ��h�w�d��wT9��+Y0�ȓqs�c)����Moؕ5���w�S}�N��
��F���US�"x��Q��r�8I�T �$�y>=��g?%���n:sp�g�*R�o��s?���A�
�d�̉8?�$o6�wŭ�'��c	�Z���-��I���]��v�����Fyr��Ǿ�I�ĺ`W�uG���;��XM�3:2��+Օ����m�#�&�c�s�~���3 9�j�H��X�k[�
P�� �<nx��[&k:�?�����_	�0N��ѡ!�'`֥���Q=ʉ���/�^��m�^uq����n�v٢�T|��A$*^�@�Y��m1H���6r	"�7��j���KlS��:r�Ko��[�a�I�޵��#i���_:.�)����Yڣ��9V�Y�.7f�W�AH�~(D�ͅ���j��l�H��D��E�mq	?�@i
���{���-���mO���z��Ѐ�]v翹^��-��x��S;�P���_u4����Yc�UZ�B���Y7Iu���x* ����e�������Q�r��hz�Y�}���e��p����S��X���m/7��z���;�����9�dΑ�8��'n <�~�_mި,V�^�lp�� ���n������%s�1�� 	W�z��1�rC��������ݖ���n�ZZ͠RG�w��v��)��d��X�sq���T�r	T�խ����︯�,�im5�s?pe��?������`�\k����B$�<U�����e\�ڼ�H.#jd��kaLw����u����c���w4��f�4r�ZJ�񉸈$q��g}v�ձ��؟������F���~�Wd�������Jƺ�����V���V�k�'Yv�
Ց�L��ecN^� I�������n*퐹�Tf�P542n)$Ӊ��X�Z�dJ�:r�b=4-�|�
�X�eY(J��JsB���/���l���/��/���|S�L��c9me������J������<��]D4�]x���n���rY}�f|Z�9t�t���̮��G(�v��߬�B��{��@!�="Ǯ�������s]X���@��p	ȱ�~UW����R�� ޱ�+V:��q�b�,�����فU�?��A�}Y�2 Y�Xˬ���ê�!dy�e�=	�ѷh�U�£�-����Z"��R��Kl8XZe��nU��%���cx|��/E}�m< h����ҙc�Tv���n�=6m�ˢ�&{�7��x��_�^r�@1|��g�٭�\\��~��o���L�3	��^�VA�w�._�o�;g�Jmc��F�m.�\*h6?��&A��*T���wU���C^�F�����P��}=	M�:�Fy` [n�Z�*f�Lwx";J��6Z���5�k�_D� >n���u>l��B	�5�.�e8x�H�}��_�9�y�]	�+�:_��7
��A<iv�)C��r�Gr#EHtQ��V�&'N,�S�Q���
�v�ӧ�F!�M��Tb�#��;ܧ��RK�oI7`�H��������ݎP�<��q��kT'�"�����`\K�����q��!P�`�gҋ=3�0��;�����[[yXJ�ɆM�&;�4n�bg�Tͽݼj[�jb	هމ�mGE��7&��M�,�ɠ���%�c�&GW��1�sg2���G�_�BxgRf�9��\�X�p����@Ʊ�Ǯ'�ոɍ������TaU����7�M/,����۸ڎL5UwҢ,���JQ�hpL����M���o��\��`�;��,��v����BU�l�+�� ��4�[�<W�I0\Q�~����E��h
�<�������HP�i��Qjn����յz�Z�*�毷"]�����'��v�'ƙn�Ma��u��:I����nt�C�)ߩv�j�YfrvW�|-	Bئ�G��X(�{�#���t��(]� �[I�����z/��r�4S�+Z���uT��n������{g��ġ��J�_�ܶ.�R�v����
pW�c�SqH�r�u�v-Һ9�\�Ǽqp�k��/��A�9��^z�1��8����:0!�����=|�_�Q�'A� �87���&)c�4v�帧/_Cl���쓖hG�.N�S�.`�����
a|[k[`���۶��
B��H�N8::�\�[C�����;��s�*��#��Z��R�c!���b�H�#�@�V��(��1�pc�m�`q��b�u�u���D]?%�����I��nz$7�T�@�"�@�U���^%_`����`=�a�ե2�o�>�e~�������U����&(q~�wpL�=Coc�1�1K��r� �$�	��2�R��������,{WQD6�SrԄ˦o�}B�U@y���W���\��5,����4�TM�6.2X��jfc�r��I�ji����<�p�\?����Zo=bK���R��D$����7�|3r�ο�;U���'W󈞄 s�5�����'��q��B��xŨC���~��~5�xHQ��П"�۴JهPJ����2�]�/)��� ��n���A�"J����Ϥ�-Y�8 ���D�)mOP5Lx�v��ݛ_5�"9��x��$1R!���2��v=$���@!���6|p�͎��e�'�ʅFP8��b:��Y��/����W5���>ȯ��=�ؕ����mrJ��*��F�1���JN9v&h�6ʃ������wNsj*�Vt ����b�e��Hͪ��!_@s�aVY�bG�����i�|e��7��9��C����cP*qq��pZ��q���\{�$�4�~�m|z��,���6T���4��F7s�=@@���d<��o�Uӕ\N��>FvO	�r�eX3{����L���b�p�2OT�Gr����������� C�Ӿ����\�{�@ˤ��.���ׄzr���W��V����f�L�BD�Hn��s���P��5�ٜ��n��+�.x�w�Y�䓼�x!����|�2���gg��m\����.(�s�S� �:��!4�Ґ_^!g�F�3ْF_��j�8��߫����-�/��|�V)ή��7�F��%�h��R��ҍ�<�)�!<� �ܚd�Đ���������d_]��;JxM=F�9!1�9n/<cƓ�It�;�J*��\πu��}��scTK��|�&��-���z�2�#ň��k�1%j��͢�Y@�@����߂����FK�l�WV����f���O��u���C���Ŭe$����Y5�M�G�>L���@'��J!@����T�]�k�l*g���
Y���o�8z���
շށ��0(���R��?���^K�4��h�M��B'G푏�T�$�.�dj~j�#sj�[��:����]H8�}z]0�-�8$���d��FǛ&I@��f��0��%�ׯ�x%>��5dG2�;ǢS��$�'1z3_|�B��ܓ����>П ������1?C����Bʝ��/�߬���^�~�%KB�O��~�l�s�*��!X�hF���e������#!�Mʟ��f\��8��M��'�x`�>����c�{�l���]��4�}�����V�K#�۾�4IV:��j ;� O�ZC�(a�ڀ�Ք3<.�˩��Ф�;�#y�^��&��K�Z�zP�]��i»��bzK4������g�^�/]/[�{*� g� ��{�d�Lz��훅 �����7�K�K�߆���X�wۯ�=�W6�K9���eL�8����%��[��u
:�<��:�l�pr��ڈZk(�}6�j�X��wN���)!7�_э�_x��m�S�F���B������b���r��:�][�H���r�m�X�%��ʹ�f�7aCE{?�P��Tz�Ф5�h
����W����������oxQ��%�N˒��}��
G�n���θ��ӷ;,B,�+��óR�E�WK��o} w%�-|����Y^5�/Du�=<�FV
T4��HUE3͉4�÷�Ni�<ۆ���ɠ�G^S��T���-G?�tQtC���K֡�7J�,F[�Z��,����'�D�}hh�0��L�8\��
�9�Y���}8���f ���ez6�(S��@��ŎOP������ҜrOö�_�%|ا	��f.�F\��d-�rI�d���FE��#8)M=�wVxq巓��2���K'�� ��m#��`�m�?�A���v{��l�Ĺ�a�S������6�b_데�W�2L"M2��J٪������sU�1�:t&��
-�=#Y���=���l4H�T��
[tF��gGu���%�D?�=Óڵsw�,
��(mDT7`��8�5[��1t{q1ݤ"�۰��E�Ֆ��Xs�R?9/�+���K��=��gpd��I_^�]ڷ�$�Wt��7�<���d*��P'��"d�YH�}!�]���F=,EV���x'jى���N��h�h�<����.q��R1��w��2P!(��D��#N�3{r���yH�9eΑ���^)h�쌔�Ѧf�:��i���%)���Q��?��� �����*���6�+��m��t�e{5v�īGE,?l}� �7�V<~; ��C�_�C+[�$j�Wc`&�I�B��rKۂ�7���]�@8�! ���C��q��"�r�Da���W\Ȫ�+��_�9��F��i�����/SH �~���U)H����a~מ�b�2��dz�~7;H�R��47�ySΎ:�5T#X�:�u� �ڇ蹥�7�g�EN�U���ө�W��wD��&�/gb�>�n�v%LLc�!��(��ܝe�����K/�h�U(��O�f�b�*����q&����.�i�ܞ�GsͰ?�3�B���}	 GI���p�f"I�|�ߙ��ee��H�|�&�	w���D����CGps樑�7ow�ִ)��вݰ4���
��k�%T�z�k�ߙ��	�	���J�9ۺ���g�4�%.M�{����b�S�ύ�0.�Q)ǹ�0�A���^
<�� 1���)�+��Z���9�s�.=9���%]��}a��P��5A�ɐ^%��4�����"yQ>���+C3!�r]#����\y3o!	�&�=I�h�A����yW�Hz�E�<�I� �8��E�b�����
�v#^� ���=����Yg�q��{�p���	�!*�ި���1�t�	U����IW|)�Hӑ�ޞHT��YՌ�'j���t�B��W��X�Z0���n����wG�V��o�/�$1a8�J�u�}$=�ټd�}V}�:��ғ�\���f���\�i:gj�v֜9��N�s��V�@[��j����,T<�D5�$����*��9��\)��6�^z!���/B~>�rC��~G�"��z�
hy�a&��;FW4d��J�Z�Ѽ�T��$;EF7@��ިX��+X*:������A%�؇)k�0�ߘ�K�u��m�/Q�d޾�߬aa֤Z&	�8�W
W3+~M9���}����Ns�'P��
Y�L��^C(��F(1����ߋٵ&�EV�m��/O���`	{����ɳ�����Ѹ�-�t�!�A�Km���?"_�N��v��X2k�=Ȍ�1IY�W�&�=�����g�^,a�)d������� �}Sh����9t��/����~��S��Vf���z*����D��ؓLX�K�Sփ.�Xw�I�u��n�_q۔W����D��Q>o�d��ϵ�גwհ�����n5��כ�ӟYz�OX��~� .'{�IX���[>��:f�����_�M���`��k΋h�׉�C�.-.y�T�_8YU0m������{yX8����Ǉ��V޷^�sDY���)�
���LP�^p�6爦�8�YM2N%��h�(g�z���<yo����ٓn�D��l�fϭ��1�Ĝ��kZ�x+5��K���T6�}Vz"6hb���ef�l�%����U�|t0�Cb�%�����yU;��[��Z9�pũZ$���aƀ�;�bIx�(�zC�)c��k����4 �1�'OvB�m���SD.�?bF���e}��YU��1������;�C��{�q���28C���(_:Jh-���G��B����yT\��H�����M�k���4&0�Զ����!��������Wc�R|@G�+u���FM����Ho���0-�ލ7\C����a:��}<�w�`A�#n�T3���dfZ7���n ��/N��:��:l�Q{�ռ+��&��"7t3>��>ڏ��F�G���n��F����'X"��Bb�$ ��$ ~׍B���W�7y�ߢŒ_ǚ^X�Xr��6�"}ńW!�W�|�l%\�oiI�nM ����q��ET�V3%=R3��4Q����մY�������9���erB�����w1Z%����;�͂�鑂��{3Z�2 P$�N�������H;l�&⎐��.�;ȝ��b�����8��Ox%#ɅPC�R��M�A^<c}�Ge�q�1���:��q�U.Ν�1��Ȣ�i�s�(���:s����G����[e�Jj����{G�0�y��Ϫ��+D��/9�cI�Û 0{  �i��(K��F���Lmg�Kj��Fܸ��/#F�
��i��	�`��T>�a��@���7kn4�d�-ss�߳-��@�m^��{[��b`]���<p�G����Ҟ�y\�Q��hUYH翖17n��T���r}a�Vo�C�*���(7�\������Yt�k��7`�D"��2������ӶNT�5�@�$�C�� �@�h���J�9�HO�P3��<�"���4�)߷X75�$`��$�c3�� �1H
�j.H��g2�6WL�V��H � ��>+V&/� 5����;�bЛ	H<ᨺ`�#��!��+�_�s;!e��PڬI��3�+wwA���h[�]�V���_Tx��W�_z+{����R��b��_����WP��T+붹9SDJ[��{"~:�k����E�+���8Eb�m�xkK5����#�?'���֍�����I�3v+Im�L���s0�D]����=��M��c�*4�;�b.��q��H�i霻�FTC��$��{l�#�z�.�k�5\).D��ԍ��<8�(U������o��i�/6�5�K�y�X�X6% ŧ��=ٍ��L�h��_��&~���Z��1�Kp��M6Hp�40R��G��֗c�g4�� ͅ�S1g0��q�'u����U[ㄻ�	��c�!��0ӭ��T|2qC��6�-Ϥ���6��5J���Cveu�׻0e�Zr��Q�FH�Y���
#�Ջ�]y�2$�'c\��[��$H�!B�ᰀ%�W\	+�����q���A��y�u�(��qZ�����A�-~���O�,�&��}��cG�''�Sd<���ʤ�QØ�0��}�X�ˁ���E�`^|�y�'M�grZX7ރ`;#\?���._�)~ӂ���(�N%j�cX\�4b��8� x�L��LⰷL$D"�����_������CI�<���rjC�&>uk����؛�(Q���~�3��\�/�K����I��1s����;Nm�d Z���2�b��ԍ��G�nk"�hJm�����$�w�ɜ�p8�N�Sp<�����	%im��P't��f!���4g~'�C ��bn�����<��)�jT=0��*����cp�)�����t��p��Ӄl��>ۢ_k=@�0O����u��Ȣ-�C�
�����n���9+	v5�Iđ�?fd�k2�y��{J�!!����
��PýZ�����Z��1�|^��L��sˆ*<��y-
1�����-����]�!�	G6���?�D�S�*u�_�&	��&�,��ئB����\rO�N��o�����&A�]̈́��uJA&�D*.C����t�2�c���M{n�־�j-è���=�f�*U�Y@Hr��C��m-HžM���)�q��*�#���c��H�|��5z��U[e����`��Dl���5"J3�)!��n�����e�m�z���iou��^L�hr����E��Q���)��BX��xzT�a��������൲17�l{���fJJ�5����F�^����z�T�Z����#��+�~vdt��o845��,_3��z�}1������j7�<]�y����>Q߈bvy�B�Y$ASk��qK_W���)��/�&%LVg��eŦD��e[��y#E���]�40�.ELz���a���)��6��,=8�.�Ӷ�g��ȱ9Rr�B�7E�\�����i>	]];���w~OpF��f���6	Ew�V�4�Z�����.o9��\�R���Ō]�&�;���ķ��Tb��izaM����^ܣ�y9��,��#U������AQ���ѐ�hx�7�������.�5��%�P���!_d�G���L:��|��5����Hs;65`��hCx��ģ�I>��IX�2�������]�a��X͜��Y_a�5z� �R��ؼ����V;L�������dܹ�+g�݄҄�tp?�c��.Z{:�aE��f�9nu����{�W9���B��BA�����N�U��~U���[�t�L���6@p̬��DtLX�D"+�{HUΕ��+�g�ҦE~+�}T	f�G]~*c�*g���(1�o��Y|���+zqԩQd�_� �J~�=�ts����0�E'h
>Y&�7݇��%3b0�稱XE��P�S��sӲ�A�����킪�<���f�b�6����!���?g�`]̧kPoMI��a��D�äFG����$��e�~U\��,��. "�k�P����+����+ǹ�����%ZJ=�q�$�s�j�t�v���_�h�`\�}N�j�X��K�/U�gk{�?a�{L���t>��1���1a%w=t+˭gW�l�^C��t�p ����.>h�
��_�2D��71L�e����z`λ����):G�T�1�,�_5���ͮ�e!����m?�(N����z��o5�T�^��PA҂�N����* �0R�Qy��  �8�ݾ�� �D�{*�s���j4��"-TkЌc��Z�"d�h0�|[��9q+��u��&�t7���Y�b�1A�����ю1­���t�8rVr��U,X�=(G�ZEy��.d�1)��~f���Q �G~E�6m�`į�m����23sq�w#��@z8�+?LRG���t,v��}y��j0Z�Rǃ�4���Ν~t������8�y�=Ip�\���(�\��[�gA`-�TJ#NS�����^���ľ#��`�����j(�,�<L �Ez���"�V��!�L�5�7�2��7��m(v=7��-(�rw~�8�t��QWa�y�!ĳ�f�R���YA0ؼgu~�����ǃ2���L��D/3��6UY����*No>U������p٩��؀;�3�x�~	���:�:2��!(��H9j'���r$'2UW�NR�\�܊b��D����j�<d�%�pm��B��X�,��~�ݫ����-�d���F_a��E��"3Cv�W&�]����*����.���|��nӢ[P�7����5s�po7�pb�|�C7q��[2�h�����]�'�1�}�6:=a�Y|Tt?��������58�t2��o�u}tͭ�e ��Oz���asٟ��rM�NA/�3t=/��de�1%��	h��ͫ��>s���}%�
JHz�NW��d����D ����A�i�MXj$4�����u��x���ք���={KUL9:v�B���:Ģ�(55�
Za��iA���?�gp���Z=���Hf՛~�� G��n��/��x���Xل2���0�j�ښ��E��<��F�Q�Hݕ�7ըL�����8�]����ٔe�b[g8ᶊ@�FP^���Y>k%i��&L�	1fbC�E4�L@wxK1{h���o�.���d�u�ku�.'�q~�"ɍ%�:�h�/��O(Jz俅-�y��~�Eew���i��〈t��@t>�:R$��������/9NFZǱO�G[!e���d�84�(�85�OLh
�k�;:x��2'$��P� o��$�\��g=/�nx���?�6��JD���^�0.��-��7 �s����a�����yq�ϓ)����S"wA����0�y�϶c�(������;�i��a)�i+mC�xv�/Q0I�Sv{:&��6<���M5��+�:�g��ȿ��(�W2�yF�Q�}/��/���|�8��}$V�e�3�l�� >څUmIw?oߐuAm���
�o�c���|(<?�� fY����~�HH���st���o2f��tA1쀟��bhZ1��
��&�	czH�c��W�"~1��$jDGST�����?�k��	�~v�ܾ�^�}�x����mCXӈX{#��f�����|/���$F�(�П���M�oȮ�����y��Zh�w���L��+c\��qZ$��RΙ�%��_0ZK+d��Bb<��֑8�=����ױ}!�_������yBG��&hP�i�X����_VՓ�EELk�R�ý�"1��b������:R����'9���8��?��wJ�b��`�f�.h
}6=�jI��I�O��2`�������^{�1�= �a\�.���I[�
���s�PK��7�W�{�2<�Y8�܉T��Lg��Cb;��?"���D��T�n��1�pP`�Z��Wl��	Z�46��s�5�wg��}.  B�����iQZC�r����~���Ք4����R�v�lC�td�sWk|�C�Q�����f#0�3 C�� ����� ��S�T�w
�ӈ%=c���u�a������YO�u=;�����,��=^�
&�4�>������?';�.��J�ĺTL�z"�\�qw�0���c��P-�e��z����q�B�0<D=߅�rOYG������c�[e�o���FQ=�N�8HoTi��d]�GH�oj��)��Ҋ}@�	Tf���D��X�R�Ǔ�&;�A����=�P5�^$ "���D��j���p�Q���aFG,к��nc�d�D\|��c�,'���iU��E"!0��
*�b����mU��'/�ϤH�}������W����)�04c��mv1�	�P�bP,�Sz �E~g���RT#Ǣ��Or4�R�� �2�Q�sEem�c�� P;�)E��� ��耑k8Q,)�~ĵ�����np绝�8�D��&`��[y'��%
�/����pb���l��UF��}��ɀ��Yv��%Bkf��ݤ7~˂���D��r.�K��3P�4����L{�v$k	{�s�r8�����Z'���G�
+mw�6'�{	�dǀ"|~ۯ�~,�|rʗ�:��W���.��?n���w�`C�3�7Pc%ȝ�ݴ�hU��g�U����<�A	��q��a��;�к%y���#�ʲ�k��}۵Ϭb+�/Xn{�SkJ�F�.{��K�愅����E�-J]~kM:��p�/?G10��~�0��d�^�`��YD£��ztZ����ǆU,,������y��
^� ��mb0f�cE�-3���fRe +���S6����a��Fm�ֱ���R�^��ׄ!�:�DJV�fө��@{:��ǉ7_SJȤ�ŕ�tRUG���l;U�:���jj��tu,�G��c�K���N���%E
�g���O��N�#��@Tk��1��P?�gy�,�Δ��(�|f�B
9eXyj ѵn�R��<7b����^]D0����O<l���}n���ǭw*��~������n>@�ٜ5���`p�BĽ�����BN�B�(+]��t��B1d�~Z1(���)��^��P�ʜ�X���oȒH����9L��g�q����Om�ζ"��N14�d��f�?�\���B�z� �1���C��u���u��"�#Cp$F)�. S+�,�֋ �
�����l�;V�T���n�C�4V�VZ��|�=�1�8a�i3�]5��n��f']���������E�1����^���y�slQ���M5�Ko#,��<k�� ͧ�WˣK-�`�3Aym�(-~�*#غh�𘭚��Q?���rč�m�nH;�w�ڜDEt{)��3D���H��i����V�@�4�M[Jz�N�뽁z��Ǫ}��E�*Ytg3#=z�z����^�/k`MӸ<�LHoIAN��j�\�ƫ��^Y͑AaJ1��<��;�l��DF�.r�ش�f �����Xm\vz����&�#�* �y�ۇȇ����vX�b����#&�bT��[���"��~�	 J�!��\�OTep}zf.���}^��My�y�T��p{;�6l(>/m{)��TU���Tb#_�� AX�9;(���-R�>A�w�f4�)�T�;�������ܥ�v���H���N?Ԋ�C�Ml] g����@ 
�������j���'E$���!X$�g���}w�t��{�����Q�X[Is�N�IEH̓�i{�lT�$�2��g��p}��ũjο�^�\б��[5EC�൪ �T!����x��X+E�n����N�h.��7�a���� �"�j4
P�7]�<	�������?��~�'iGG�0�1sw����Eq���O���x����=���^iN���<�(�ܮ~�4M�[.ҝ{�Gh:���"8E���V&H9T�ݖ/�[Ӏ��:^ۥRfh��WS>B�N���Nr�	n�Qd�*��#��P�ߒ�@�7��������i�y��++Z�ZV� *�������%�s�����n�u]�;�Y�Z+y�*�gI*aݶ�#m��Š�����^ڢg�0���qebg��@����a�%��*Yd�*���� �G@�g�y���� �>B={�5b�}�&7��5n�Xd�aaU��8�	g�A����|����o��+���b���K��Z���bw�*8B�U왏�@�SPqY�:����60'�/pؔwsf���D�;��.���9�U��/��ґI��o�;�6f�4~�w_������j[�4��|��Y݋	���p�7���a����߹�$����p�b��bZ��	����v�`�w?��a��11�CscӰ���kȈ����{���RT���6E(z=X���Rn �XC��~��a�'��Zk��3z)��%���#y��\��eN*�/�5�����u:KWG���=�G�h�v��4�^3�п��m�+�Z 𡵢��>��{c|�7x"�WO��v�	��U�[�؏➡��S��|�@l�ߙ�@�0c��?��V�_����N��T����t�3'�H�g8-�9
*v��}��׌sۧ+^����Q�7��޴����E;H����FHh�ۡn����vv��Di�y�X*��f�)��#�w��펨�r��gq=@�e�ݢ �Y&�h�ӵ@��`O�*�<U;����?���� ޙ���hYi(����2�qO �S0�)U��I�Sh�F�g�3!��74�G���J��?��"��͢>HVuK�<��%���7�q����o76u�2ͅd2{��y]l"���|�M��mZ֗�I���%���#�t�cH�Ѧ�n����B�`P�* e��~�D�d7��­�}8Jc���`*)��/� U;sQL�ă�Z�-kN���i��zPG�7����g>�4c`��
o�t1�84	�4J�_��ul��5�w���}H�����PL�|.�gɴ_<��	]�@��LȌ����|؊*���Ǝr`�����e ��"��&�*�.��ִ�����R��@�k Q�S6N���V<S׸�f��IkEG��Gm���>��5vM�A�a"��ŉ�k8r9c���k�G^(C!#9��x��X���&`SU�-�0�l�(���_�U�-��p�m�rU2>L�֢pYԟ�����(T��7�9�8�mbz�;���.F�C0�@'#Z�8$���g'i�903_/8��i���aO���b�����,5D=- �\��ׄ7Gx���X3'G��M�3�淲�E�!�߃-�4����ȟا��H�oF�Yu�V��Jxs�A��p{�4�<�Rs`f����ɢ�+�@�g�M}�p[.��{`��@��Q�^���;�)��l�yQ���X�0r-Մȍ��<Evt�ɡrzN[�|G�����AB����f �����H*��qs���	f�IHe�1������:pТ��wV3��Զ2���M�(��[�M��O!g��처C^n���y�����N�h*�	;��odE��F�- KN�j����CWߜ5�B�x¡@�6�7P�;�(2���t�'"�n�nO��5Ey0}M��[3�"l)�0w���#I~����>��(uAS���/�r҃�? �����L*�ه��n���ւ��,6W!b�l�KpG��N����X]�D��)3=�`է����`Utt7�df�灱�v�%tP�
і�*p(T�۬Jg�УS�����j+�,�A�x�Zh�Z`���|�ޭ �}�
Nd���Z�\ ���) �&
����
�>+7N8�Y��I�F@���D����xp*���,d! �հ�P��������y��N��sƯ"���ؐ2��w���.��x�
i�W��ѓ��=���sYrz��ն��x��h)x5gD����������N���FM0��(��xRgE��OͶl&��.t��_ o�߳�b�3��/�\���6�br#� �N&-�h�+�"q�*8r42��z2�A��/��Âv�^<`#i����� �ub�ޔV�񔠈
(��I��P�f,�u�"��s2e��UO�q���o�=ѿ�DtQX�	�+Ž���?Šкz��b�/�Pf�������'L������i[~��*��2q<�0�:��a��J�
w�� F������b���vm�6�	
�r|��t��d��J�f����W��ރ�4�o�'R���Yg�Uu�:���������0�z���\�	ʑ��D7����e3����0OC�ԥ(�)M&�7��E���E�%�H��#��ڹ!�1f>�\p����~�T4/aPoQ����=,��vj(N�%�c�34s9�8�� ��tP7�~��3շ��9\��ى�rs>�@��Z;��ӌ�A/���Q���o�ǃ<<C�9�2�`~N~|E!��'���<�g�y���k:侴mo�V*Vx#e�c��7���>��Ъ���?��^�nCQ��!����}b5�xMŰ��9?y�K܌�g�Cz�'Pgo{ɢ[��^��ރ�-���	��!KU}Ħ�:�b5��a/�k� ��O@
.���em}$Նu��ɗ������&�k�IL�`
Ɠ��Ɵ%(�m�og��Zn�^�c�������TFi�c��BgQ�S40�R��s�%��֩�ݧ5��V=��&��l����&u�rn�Ұ���a*~��P��L��c0�9w�7���}�۩s?�I��}�y�
岸��ݧ������"Bu��lkK�ȵO��D˯m��7�����	l.�8"`�-�\y��B	��4
��Y��s@�����%C�d��yX�G8���{U'�t,�WJ��$��A������o`3=��=�.WޤߧmX�h��
�Ī��
,�bz�\�T
���
H����3���w��o��)Ԥ=Ř�����bܢ(��p�A���m�D���Bs'�; ���3h���w��2m-�&�/�'�[�aAPIx�Z�O� �~��6��`�� �d ����I섻#=E��D����:#M�s��!6�_���A۪f-\�s�t�vO�Tw��Gb2u�Э�O���+�j��e:�``(�,��-�-kv� �#�hv���<\�_J?�oξPM�U�|�B��J��dp�.�>@K7�,��>F�F�,�8^�.�$ޏ��lm��3(E���>L%,�kM�uzu�Ns��ne�+pY�d�{uw��*�HQ�Koi�a2�%_���;ԶY`g� \�.e:��I�2��rF�@@��T�p�}�N�J�in���.��l�IL�GUKER]�-����Xm��;���!��6���-ðz�����_��p��~j#��2������$��7�7��&�4��>3L��I	L��T��p��5�\7��� \�궖Z�FDiౙP�H���.#�3�UX�>���ǭ�[�g7<�N�b�����SxK8?j��`��իp�;r~�׷���|BA�Gp�q?��"<����
� �3�6�Ķa諯�q�ۉ�XA3m^Lv������2��VM��`kT�x1]\@!dQ��joJ��J~~�w6ȝ���~��3�U��a��,�į�Vxt5�]�OrM]��q	3��%nHr�*�H$B�l�]{x� �Y}�
S�j#����1Z�p�L�����z�mH�� ��wW�}0�����ܾƢ�bLt�@��,F>�N7-��ʖ�wa>�j��M�q]<�H��U%�,[E|)֋fjCl�9���p���ž@y�uiJ�fO�Qr���϶��[�!��h���f���#�Qg���JH�J��4E*�{�\y��	Ţ���45�nt���w�~�������\���'qDM�xP�B��Y2+KS��'�ӆ�Ķ~D�$�r?[�9��~��OI`�Y�Umԉ�!�r�T����8XN~��x�/o��H�*�(ƒ�VGE�0�������eu�M ����U�K ���A���	>��df#2�b��Hu����Z�jS�PZd��ڔ�'��D,�n���u�:��T��G��CvrM��g��'�%��/���WM+*�Y=y{�f��0�H�O���m���NՏ�bs �H���Hb	��Vg���u�������4��|v
~
_=;`���F(0`��=潨J�|^h���qV���@x.&��0�y����_�[ZP���V�'�M+�%��dO�?ڣd[�L��������a���z�����@�M���l/�h�u� 0�W\k;PtF >p�-�k��$y�Вe+����h6�ЭCc�R[o���״�j6!��H��}!r�1x�V���_�sq������<�;P������K���.��d-���8.�PP��Д�Э�ݫ�,�l�JGJ�A��N��;��:O	r׌iD���q5:z�.��j��������>b���d��P�.�Md�ʼE8�=9றQ0��z����Jq�O%��Ȥy�$���g�I�B�!l�?�U�JTw̖t��hV]�9]�r�\L,�|�ֳ�Rs�<1_ݤ�u#�y*�;��92{�1���^S��Q:Ha�3�'�I�� ۃAz,�j��>9j�*$՛�S1ZZz�N��43af��ex&�&
��(���D't�MJ�՚�[��M��) �Z���˂��W�U��6�?� ��(�d�ʝR��n�7/���Η2! qPR|n�'"��	m�F{='el�^�Ŷ���$.5�����RJ�LF�z9�_9�
�1��JRH�d!+J$��q�4^�ƥM�`���a����8�쩼@�-gk a�Jh����!v�ـ��S��G�OI���!/�|S|e��WK�
Z�f��=&J�!1��G4N��ަ-�;ﬨ�t�,�D��p6!�w��N�|$��<kb#��� M��2]G�l)<�o���d̒����|����zr\����i�p�Q��wmc�ǜ��uCH�`4x�jDِѓ?��z���5�?l�y:B�*����\LKԁhd���G�1Ƴ�����3���n�G8tNZ��F����`�~�:6�zq��ꏙ��1�^K��a)���A��<c��=<q�~(I���r����
��sg����v���;����_,q�r��Pv�}���LiTO�CQ7��7Yq|�z�q��@�uo�ȵ� ��*]��O��5'�$*��V3+Nf\��$���}�}��kD���(S(E�NFu��,Ĺ�}M��{�Vm�.��2�J�?��l��S`���-�t���j��;#	���h��D���#�������r"A��$��h��o,�-dO#�M��9�s�8��<̈́��Lz?˹l3����q���8�}�+����$ ��������nK�T֕kȱqa&.	�#�3���,�����"��Kc��p�_.ַ���`2�r]�!����똻��x�.�-�n��<�z�B���֙���<`>S�����}lR�����(i��*sZ�M1�[����8xG��YB8w��S�%Fm7T�no	?쿲,�A��s��w��Vߔ��a+��X5�(���ZPl:���+en���n\��-����L��3�55 }��e�{I�$a�nm�~©ʙ6���]��w��{���E�D K����Չ�n��(Iy	߀c̝�V�F����@~�	3��|�"�Z�W �
�ѻ�
���$r�~>,Y��@␪�Nz�(��H�Ӊ/����T���[�����z]�H�A6��O�)gx�fGѾL�2��ÓA��㙧�rT��͑s�0�����9xJc���F�E[�� ��?M]w�[��H��=����z�XI����|�ٴ�gM�:���׵,���B���@��Y-si�u����[*\��?��vї�n��e�~=�J�V|���f���^`�DI}�,�\���+��kU䆪� ��B��N��:�C��z]o���A�#�I���iB�U�4�%7��k�l�9�W\�:R
#���)�"�Ya���̙0�s f�Y�%Dk�	�Պu����清��/w#y]�,⿄��Un����)@;����̔�W$^U�k;��nLkX{b�����ɢ�an�����8���o~� ��ڑ�L0��ݭ��`��.1M?�>���b�M�|�0����\�s�U7q����f�5g��F9��;��:��|C�2�,\c��`j�)�۱\FX�~�3;�~"q�mB�1s�4�䄎yU�FI�Yl�������1��0���`�w��Zt�1HO����A�s�Kb%]�ץ/K�^$0���h�+<|�蜔�Ha�V`���ɃX4
mf�]�,ؘ�w$YvRJ��9bgLŐw+/}��a mLj_�PT�dҝߕIl�n�*S�&�d���F~�u���S�E��D��zͷOm�<�d	H��t(�#>Vbߒ��͚����jbwh�u���Ʒs�s,�X��Fӵ-| �PȉUI���_��:Y�8�F�VR��a�
�.��O��g�X�5�j�[�f�o���ϫNx%ػ��C�L�z�X��V��:_��0Q[Ŝ��R����0|g�-��� Sq-�d�d�S�w$����x�t�Ѭ���)�ȺbK:nEPI�|�_RW�
�q�j���2�À�����$L�)#5�/v�f���r'~����8��Fc��?���S�o�l�bWgx�p*�L��𷟞��"Y�����@V�7��:U#��S<g
���	'F�;nFh������(N���m���k]	t�FJ�E�FH�3k�����Mw�&���ʉƭ�l����<׾K��`�ٯ�Aˬ��2|�_B���3���w�!�ߕ~Kb!�M�I�$Ĺ����xF�P���Cޱ� ����s�)C�{�	20�!gdX56�9�y@���G��1�ݕ��q�B�1a"�i<`+�Z���d�,`�7����4f�@��Y-���>4�$��kf\��$��'O�]M�|��M��!| ���&�L�-u&��),2!+��Qsg���C�Z!Bk�A"֡e���]�}�.�����B����x�6�1
�aX�`x��_i�J��Z-Z���ݢJ��fԨ��Z�(�V��;(�'��.20q�w��z*0���ནX4�ۨ�C��A�W3Z�~��J���2G*�:��_�]�<~
�>9F pb���bGC�1H��,�um�tQ5�.�
�'��7�sS���2�/Ր�@
�9��'Zb�K�$�|�N�&QhRxH�Ӯ6����{�Y��#eO�CqX}(������������|nY1p{G]	X�i�����=�{)9�O�o���L=h��{a�ʟw8�����L�a��W��*���n�o%>���$�E��;*;*m9Iڝ�Y-VFQt��p0�D� DB�����tWW�[""�\%)8�#����I�5�I��׏�c�E��O��\��J�P�T]�]�ԓa�j.�f��2暲��>I��U�<+���`l�?�Ͽ��VQ:^�Y��7�t���D?���#N|̳�3V���nG��4qz�s2^�a1���9ѿ��<>��k��w�b���o9�"��7~��(�K�<�b��!�M70�JU�ٴm�����Pd"�ĝ���[�c��f�'��Z9b�h���
��w[]��C�>#˧�c����&0YǲW�oޭE�%8Î:�
�Jd�4�|����x5�}��/it?ku��?y����w��B���G��^)褷�5$��ucs�@=q5n���5���Ø�<��St���|h��J՛p|�R�.�W�W5��/�QY�I���'L�����r�G;��A5�K!�kC@b2�w�mfn�(�|_u���)��$�5���#~�y{�Ei3 �w�-âR���j �T�U%]��'��t��aĊnu4����G�7������fJ��eB�P�y�h����F��\i8Irp(�P��h.�Bej�?��g�-���I���d�"9T*S�M@�@�+���Y�ϟ%���͔M]�sdߍ��Gbq�@���3Ωa{��~+�޲x�Z �[QD�FZ��[4(�G1D֋~^�7�ۀA��'qMb�+ߖR����������4{j/�-�؏A�ѷWt9�}���=�����T[,"�U���LID�& ���N��$�#��@,V��]�?�Rjb��G��;��@���)/@0�3`���.x$�ȉ^�(�H��u�Dh�R�ͽ�e��������p�C��h����Y��ȕ����:Vևۤ��A��f�A��@���Uǿ6!jԔ�?��\�V����^O.�g����)(E�"nm5�n���#R��9����W�,U�䔳-��Y����r�<��(�m^x=;(�=�҃u���q`�˻Fj���\��l05��{���(c/
!�W��h^��@�|K����%����bXMi��j�
�S�����|�%_�!����}��l
'6� 7����+-�|������@���]uk�����5���Ж-�4!o�0$i�_E
w�0Έ��6,����;]9�j�N.Fe�!���"�h氯��F�?��.����w��D�]�����aj7�qj����$��
�q-�i���,-�?W3B[]G�����Ԛ��
� ���1b���֔��Z�T8U"Ue��`����>n�Aï:�7�<��Sw��Q�<	_��hL3�ǛS]�ynϚo�>$�s6�(�pL�7"b`2�
ъ�/��'��xwd�\9�=l�5�</q	��D�M�u4:B@���$E�e��X��a).%(�=�Y(}��ř�D�J�W���G��Q%�Tt��EX'�;~gM��;iw�s)՞{�<.f~Qnla�㔝n� ��u���_0t7��b����F��̡;��r[(GL!ͩf�E�p/���N����S<��Fl��vJ��j>�Wi��d��D_��x��\�o���2�+�䝸�O�Vp\����΀��+���Q5��� e
��MH�- ��r�2N�۸��2�� (��f�)rAHM�\���@�2��J$�� #��&���v
8�*���D�Q@ܳ���<�V��ޙ�*�@����-Ϧi�cK0z�_:;6�j:�vˬ�oͫ@���s.&ŋm���D3N�����Sm'),�s\ݤ�<ʅ�ʔ�&�͢�i�.O�D�1>l;��˯s5XU���T�2T��Q35L�%�f����ԡ=f���f�aXJjs�[/����m�`!���wۯ����NQ�H��X,�0���ˡY���|$x~BP�����O�6�ݚ�O@�0���$ܠ�],��0��G��U��8��~P������)�pC�����*�q��7��$*ׇ@"�P�g��Hw����""�Y������g�9�%�k&�����)�3A�$hDP=<�NF�����u������L2ZP>e$�yFPQ�K��3���Ǎ�Yx`�#ȴ�"1��jvˊe�`�$KdJ����!+.�^��o�EF��#H�ye�+{a6H_�����'�I�&ګ4�c�=#�d �{5��o< 2D��r4 [���C�-#"��Vl$�45"�"#���Y��U�F������a��=6=�Z�te��Gh����7=h1���.�ss&��f(���#�tF��B��Q�	�FSu�`Z>��L�����]أr}�j�p�f:"h��ی r�O#��q�j�~�J{
rcè�Xq.&&����!$�����A�خ��S�ͫ9�'�L; �;��s�w%� ���[g�5�e�?z_k��̎����U~�ȺԚ�)��������6�PvsJ@��2֜hY(!�Д�����у��@��C`��n� �2�*0�0�&Ē��$��!Б�F�$>�Oc�8��==(H_q�U(G+�B4U��L9��@��6������z8�x�MECuA�s�y�*�Eh{�|�Ϳ�V�Nk�[���/k�U�ƿ
���G�U?�e�9�d)h*5�(� ���������F�ݏD�y �n=J~��0��F���D�|����d�H���^���q�`X�";!�i�Sp�z�����<=��k����
_�\/Zk\q��`��ӞW�;�R0x�����g���=1v�_�!�ɶ�C)O���xi���/h�O�����XoM�����W�:#cZV2?(�E���VŅF�h��p��7!+�����4���O��12�zn����"}���r��J}��㕻]���
���7}1�>�Fq|�.�S�r���'�i"�6�Ό�򭷺o*V�H����ټ>�HE����#����|n�S��ޮ�E���G��ڇ�ꖋֿJڊ�d���3�zEc�dgv8A6�.T)j���:"ݞ��t%4�o�g� "N�z��ڲ+����6���&+�3���<�`�@a�!!��uc0_H莴�c?�b������ɞ�>l�9Fj�;�T��i8N2\���FP��a%Rvp9�����WfW��7hf��o��OG��<�L2�zso8v���>4J0��Ϊ[J�[k3�^a���6���$���ڊ�e���8�"�?p[g@�v4�������C_a�gN���L>����+�$b���;"�+���-�0�Ѧ��]�d����c���W�/*^g�@6�XÃ�&[�������0����j9�^o�������A�Iݕ)�Y����#eS�b�8;2*0.��>H�FW���z+9n�12]���)�5�v�����pt.��KBGih�����[�ջ�mJ��=�I��^|� }����㿊�X\n�9i��cs��k�:���u�����.#����C@�?� �Ŗ%s�hb
�S�l���I�x�{1��l���1:�Y*�=��14'[4ey�G���B��+�m��!�!��H�P�	Z:�fD����D�g���J����\�XWw��*aQy_D����� D�N@�}�K]�������<�QS�,�����aP�G*�=y~k�mZ!%�6��Ý>�r�%�w�!t���WһB�X���������l��
�+��o��2���T�?wX���S#�q�>��ce��
�o�h�C���`�=�r6'��ں�Yq*��2[����W�→�� ��|m���Jv]$h���L����㖊���H{4XU5f^i�BC�!6�W�R��80 �$3��x�<� ���-�O[SC�n���H6���.�����6/�,!6�hX���nC�%���3����.��{�@Jr� ��E�@;H)N�Ԍ&��c��j`+z[��̥u�=���(>pL����^��ht}�)n$@\SP\�:�X�X�r����y'�� ڈT$�Qd�;:��G�
�f�q��g�����/�l�˿��[��F�e��ʃ��%۾�0�:$
�
�"�8T�U��(�}��gF
3��.:�w>�I����Dc�A=�AaȞt^S�H���E�el��LRx1��z�TN�������c�D����+�:ꮗ�K1$TZ��Cǳm����F��.E+Iܦ���ෂ?/p`��g'B�m�A��=�����1QM0�~�����Y0�zҺ��jP��4������(�.7��xu��Ԑ[-+�?F��8T$��B���f6L�%�&e��Y�6� ��N�v�'?Lc�����q��c\���͞>�ס�F�V�(�BW0�F�Izct�=�����xn�����k��O���j�8nu:�d�w��^ |�����g+��0����RD3CsZ��ʆ'��4�$�e��
��*�x�j_�ߋֆ�Gn��Jȇ��C�6���^h�g���̑�1m�8 !���G�B%^V�M��oxCXOj`o���M�3�f-X�Y�.���S*{ye��I_�eg���?^,Ycu1�)λ��0����bG7I��[�� x�A�WT��,Q��M_Ңp!��K+�������j
�FN�!|B��c���l���mg��,gxb��I��>4�f�(SC�K`���չK�ҷp�D� ���I�x%��4���3��%���	���S��t��r�G7J�D��~ �*1�o���HDM\�g��t �ekCQxPk,%o���	7���_d�(e�)���`��1���x��gV���;i�x�_٩�E�^ޜ��z8��|�Е���X�$,��
<ں)�b1�2ݟ[��:�.C�	���@;� -�K�C��p���&4wnNΪӀTj-��b��h�����i�Lv���p(��Ɯ��)�mr��ѧ<��Y�����B�x@�T�UK'�n����|��!Ԅ
�=� �B��A�|W�}�ׯVI���j�z�{S�t�jò�v���s�q���8��?���������0�R�o1�m���R��~��9n^�nu�J���F�s��v���>�����fKZ�3�'��N��"*"�5,a�^!]�P��d�^�?Xx�r�7���E=��m9�epDPI �gD�b,I���"�D��.	����� Z3�p{��z���Vh)#��)ږh3R����T��/%Ҁ��;��KO��
Ѭ��>�Jd[����֤F]�)0"oU�Oz�d���ڄ�%Yk�:2��E����ڴ@ͻ&Z��* ƥ��\�{���e��^8��sn����&��o��̝}T�%���f��sY�{���Ki�L�-$�6z^�w�O��u$�9���o'��$���	�1��V�C�s�}��5�R�o�_�HO��7�y6
g���X�����g����Y����gHqN<�d[ c�ذ����~�<Or��	E�ߠa	*���ݼ$,�}��`�ѫ��ݠj�f/B�g=L���z��*��N3_%���\_d�z�Ƀ*��)�5�U���{�:td<���=X_��_�M�>��Y`�+�F0ֲ����[�),���:5'���B9�#E�|��ǽ�ӜX���?����0=
����������r9�}��d��+n���k�z�I�VHU��S��V{T��i~OC?i�@&���L��S��e{��Ig��S�ҒqZ���#
����<)5��xQ�VHV�'���U�:l�j���y暣U ��~��߆���B���}�/����Z��9�U�����mD� �Ex�˸u�̞i�8��=*�B��>e�uz�v�F����z��O��5�3�0wV����d7�^��/U�4��������12l�7������B\�y���+��1?�ѥLp9I������`��G��U�D��<W�F��Wu�kk���9|UX�^AuD-�췓��94ʥ�(�[�!��L�m`AJ��H�L�e���X;Ǯ��M�	�f	[���l/W$���'�*w-}����~��,��Z�'�3@Z���	��(*�#����L�j}|q<�?��8�i�k�?��Dk�h��:�TW_�D0�v��$�hǆ� 9��������@u6i�HE8c��.!�VD�:����f�f-@�?�&�2w��4$�=ˌ��PA�������_�N���b��O<��G7oU<6=8� N��w���� ����~G���UlY�b�`Ĭ+#��K`�P�/�0�t2��	,brm_zhAսfa����u�v�������]�nQkQ����:��5�J7�5|�/O�h>p��,XT��M/���u=�zV�V����b(٤Kx��1��/׌�>ȯ;��K�,���O�>�S6j�fXG;L��/J�����Hm Ĺ�ߚx'���`�U���/�$��a�9~+A��;������0��Gt�	���K�us�<�`�Ar�H>�>�<��?�/󟑶����cŖ
�8��~L�8bPZ�ê=�߽h���k�mL}B"������]�4�gY{ڂ��j�p�E����3�gpATM,h�/�*շ�}d���R0(��y	BL�{�M�`��;��K��
Qˣb���0���`5��ϔz�`�6tI��̯�=�˂n��@��4��l�Șj��рy����<CA2Y��O�7h
�b�X�	�������t:�5 }�xj:�nw��2Z&1^<MS�N�O�_nH�����ץgS���EJ~��0����������ׄ`��&Y����o%+�H��%��\M�,e�6IG�h3�X���:c��cX��+�0�⸀�<,CM��?�⼗*����ZoJ��'����C2D�qk��NI-��
���;	�u�5w��^W�{Jg����Ȣza�6��	��0�/;Q@��<U�����7n�k��8_�Z�3���lmb��Ue5kg D�+'"�Ո>�Q+�;��O	4h�4�O�e�N��ݢ��P.J���@ͱ��'tZ�i`Xy���VV�A	�>@��ںi����8/�����]{��5X��h!8Y��U���q��h\	��jqp%"z�4K��ss$�@8M4�QG���!��ྦྷ!�4�,o���+���v-�{6�=3�9��L������$j�S�=�G�L�_c����n�1���ʹ��Z��B�b���(gᎡ�����k�)E��ٵ�,@���C�ֶ�b��X�%�I�M1x֗��/8�|�/�ؼ�ՎH������w��z'(�xtx�L�aC�~zJ��ݯ�A��KZ�l��Ҹd�[F0���'{�ms�'�*9���^��g2�oJt����"xWgs�?�=0��m�����9�X�\\0�N��-	1�&~�tKѡ׏�gn�I$3U�+ح�7� �?mq٢D��iN]�$��i�@+��B�H�Fӑ}�n,Q�뉒��r�A<��h�u��%E�)ȧ����yT#W��Ⱥ���N�,�<k�x��p�A�G�}�A�����yi��v2���Gp�P/����0��.Gْ}�h-�czV���v*�QAb���HA�!�V��tk+N�O�a>����s:�I�n���F����\�#�s��*���I�²�����E�-j0Ar�	WF�ދ ��82"��A�wX0�/S/s;�8�ϳ��tXN�ӗw��6�Vz�a�U-t�6"�������S*�E�_���f����M�w�(�m�cݶ��o�1����|�i���5��8�T�U�2��|P,a]�YF��y㩀��"��
{����Ʃ9�J�����/��2���ձt8��xk����ve���w��G�̏���r�Ԁ�	~"7��<APz�dX��廝��T����/�-��Y����!��c����G;��Uy�H��7��\Q��7��[CF���|�R):�)(0�� {#������hEyPh���R�H�+ҿԊt�DLl|�畕��A��W&�X�R�-�=�.q�c��:'B0k��"��n�R�*�&���y�|�!��MyfZR�l��O��}���(��P��A��/V�q+d��yi�[L3�ܰB��re����Ei�lV���^��������Z�@]��eV�/^����c1G��,�w�-FN��EDc5x�h��C�Y=y|����gd}�M*mr�E{E4���e���`c$�?��$`�g'4׷)��߄��Ծ�3��z,4���u���s�<�Or*\�կ����fL�j�C��*5(�z�xK .Rڬ��pȳ3!�%��:�<��	�1P�}i�u@W�W�݂Z;�lþ����ڬ�<ͨ�|��9���=�Pn����g��@ς=�_�t��G;����˙b o'�x�`�`f:��]|�"���v".����QF] !�ɷE,{[����c&������I$N3��2Z���*��*0D,���ײ�i]?   �}���s�ѵ��$s��<e�9����4V|(�k᜽�z����X�b<�^�rKǧ�<
�(���#����t<��7�Zȭ���x2��}U�1�c�����F�׹�H� 2[��������3m_�;��
64�� x�^�l]�c��T��ǟ�ٱ���f�L�������N^�v�v�:{ќ���FH�������$0�ו!�@� U(�H�!Y�$&��y>K`5�K\&�\ޥ �~�o+|v����!��F�Hfh�0D���`�xG�4�{וl�(�n'��
x�Ƶѯ$�	�$3�8������s�"��^���7%ͨ����E���ߏr�{��R�\�K8?y�Z�6S��ռR�3�ל���~��I�9��X�N���0 ��M�BX���f̓F��R����g�̸�$iI��#ٹk���۲ʅ�1��&DzN��E"���@��Ѕa�@�tr�u��/o)�H��r��R� ���=M�� �����G�̞Fav��&u#��G`g�`:�UE��.��.��
p?������7���zEY���W����[k�9n��) q�I������٨:�K�)[��IE�tg!�t ����"w������t8p����)�Qs�W�� �����j5{?�Cdgx&ˊ0��B��_҄a��s��\}��On-�VDW\{��W�ā!p��D"�A�:��i�O�q�B������=U-XGP	�K��X��a��uD"�wL�MHz��tj��;n({NY�eQ9f�W���\Y�Q>��_#�'�;?4[�����vЄۺ�RW��dj�l������1�B��O	Sd��(ꟑ\��Kdύ� szX�w�7Ԃ��4M6�BXlf�}�/!��L�tҺ��J8�Y��Y��NX���+�g�^�yL����K!*�b���֋�Ԑ	B7�N-i��p����_J|��K���g+IA'�>�0��4'�3�.��v�ݒV���w�U��9<����)�w�g�M u��3R�B����}O�nQ�AX�ݶ�P��S��
|��=	c���7�Q'}s�gR�{% ��� r�/��:҂_Y�J�	��L�m���CM�K������O��}��5�/W��2�+_qi�\JB�X��`�6��|���o�2������<��B�Ќ$˵pD"�xG��u�ЊL~ͦ�4�.d�~���ǲ
���P� Ֆ�1�x�=��?�:��'2��ߝ���E�P0f3h!�Y��32�+����>o.����m=Or߼гg�#Iy%W��%��O�PIg�A�����.!Dذ�$��/,=�3����;����c�6����C��09�[�H�e�!�Z?5��g39������T�UQgmOՇ���h���aj{9���b��g��C�imt�`|:�� �������s�f���5�:��֘3݋$ph��]n�[�P�8Ĉ�5��t�{�wsC�C�=��,�����ۗR��6�넠�~��3Kg��~N�(��r3�iu�m�)�u֊\�ԫ[����cOj��hE��D˵����^�(�.�bA!���!ߪ�1a��4�N�n�<c;�����p}M�u�^�U�ڑ�����MYs�.��܆��^����YN|�+�5<T���q):n�,�N�wr:�hܯ�P����N�r�6�t�M�|�QQ��O��fu���o�%z��x�����nr�5]����j�-j�j̚�x�J���!�^��刋�kMTj�zZV���!Y��-�c���i6�������<E$�(%{@[���
q�2���%h�;4Ld�H��ĉ��Ş��"B��@ط";>�A�и�����	;yVbǋ/��G���3��+MF7�%ˢ������*�ek�#�T��c�s� �]�[��W��{�nN ��\���R�7T[L��3b`�q�	���i	Y�h}���H&��k�9B��4�5O�<�����Ϛ�/�b8�ݖGq%����Sب\9@��N��7J��#�1��	7{��&]c�p:h��B�}9 ����Brta��F?r��^Lm��8e���Y�"�/QZ���i�=P,<%�N�L_V^�H�@�	K[T��XauHpn䚔��[������RhN^�vE�j�s��٨v֩\A�'�;�D���t��)We����Wl�3m��5?X��mD��!�������O$�Cc�օl�L{XǾ�i\�zh.ϳ����z�`�2�D��祼=B���s�-��O��@, �}O�R���"f�*]nW�r��)��&�.��:S5�l&8����_�!v�o��W� ��t�P6<BK>��m��Wu6R������٣r'b�{Ǐ��cϭ���o��q��r*���o�58!��-��{"��tr��k����S�g7bϬ���X�Vd�Ɩ�v��3�˕»��c
2��t/��K���L��>�C�H]�R�5��|����b�L�҈�r�*S�np��	'�Q���z4�ny�k�[}<���:�K{T�x6��$�;VG�����4R�A�	D�H#��g�	!\��̻�'�ʮ���1l�z 9���U�f�k\;�صV���t���`���j�����m�Y6o�{��!i��>S��}�ڡ
k �K����_8�cr�˛����הM鲍���y~sV�z��:��mI��l;0!g[ޖ}�����sQ��F~��� �U�<!�=��{M��V� ���B�1������~��e��JTeO߽iՖ�(�a�x�B�nj��[e��H8���ŋ[;Dc{k񔈳	��"�l�ƣ�,�;��C34~R�xnO
	z#���a����8g X4}"
W8ᚭ�ͧ>#G��������J���������O�v�I��oѶ�J�c��vh\(���+�1!ܺ��P�_ef6��Bx�f3���^��EJ�|�ٮ;��e)�X�{p�|����G��Ӄ�K��(�*|ي���ˈ�|���(�s�c1g�ɍ/cGǖ	5�'4��T{a�1��X�'/�:w��- �]���/j�+@~<������ʗ�ݶ�\Q���c�^�{�D� H�s��D�2YWsi*Wf��rh�I�CM/�	F�:2P
�G�� p�&�H����?�!�ؕ��<-�ื��W�V��3x�^ָ���~ߺ�ٷ}d��l&2ʲw��Eй������#�^�.-Y�ຏY�G�?ߩ�O] �rv�*f�u���s���K�S�k�����<�@�i+���;�_�E����E����{Ƙ�G!2��s^n��B���#-|�;ɹ�Y�4�}�5�g�j��p��i��V����2�>ܠ��g�w*95%��q6�$.�y������"H<�"�x�ʜ�e�ڋY����W�um�:����-֝:�')����egUћ����ˢݼ��+b/����5���,bt����
?v�o����1x��.U>9�P��	�n�Jߚ�I����i�5[!�r�N�n)d�w'��
��KYkkB�r���	6�9~rѷ���]L��hw�p Ʀ��(M�if�i���8^V��6��3�7Ja�r��c,sݵD�k)��+G����:����:�Ȗ����/"*���V �$��#�PT�m�?����s1�~j�f�	�����49Q�CЭ��t�V�C�vtLUsk_[~�ZS���P��U�Pg�����9����I��{Ö0@�\�.�d/уG�v��B~M�j��i(D����ue|�ݽM1�MT<�y�]O�*�<Q�����k�Z��ZJ^�a1���vDXu��@���:����&ttه� ��#LW�"~��,�![s.�2���x9�-p>/4[X4Ԗ�O�c��ǐF(��������0L@oH1�\�vw�v�����b\���)h���0ht�d%��#�,�[�=����l���6g+�	����V���ֳe���F�G	�i#�� �~��k�ɓ�m���06zy���������9%��]՗���$��S?#�>l'��ڌ]� �b�E�9��S���g��$�d�����u�(?c@��%u��Ӑ�~by}�P@G���-!�j�5`)Ƶ�@$T�n|�񥊛�5�6���@	e3���=��.�'����j�?ܬ�_р�,�ןY��'AhOu�@�,�Q|s�@|m&���'��n>��٨�.q�D�r�����3��ɸ�}�$�?r4�^~�5,���-A#��l�"TIa0w �g锄:��:���Cp����.�3��;kw!���L��W'��W�ը�@�+�k+���CĲtm���zʦ����(%�����̵v(7���RL�&�R�奡5~c Ӥ���n��:%�c!$�v����(�W������Ng�,������$!��kw���7����$<��R�3Ӆs�%��?0�
b����	�$�����lU����#��2�QjA%�Z���쩗�I���</���!)Hi���4�^���(�����B���IGO�i�lcUS[j|ۂ�[��s��ra5��`�\�5i� j���	�t]�lq�u	�{�F��f���[nI�:��{ꊬ�8Q��S���t�c���V��PuV=�������o�I�-B�I�7��6?A�GZJ�e�)
��JbUa6�44a@���p�/r/]d��x�~UN4�KI��G3�w��f�8	6�"���.����mL��ˬo�.�v�2@6Y����!���őBo�mc�]�8�C���4���y77�eN�?y�N�\�/X�p�,d�Vw���9�VV���1�t�ǹ�rL>$��Sfuc��@䶂���� �:�	�*�7Х�%�8���^�dyc�-�7�����g36uc�uo���a���v�uf�J%U�3�����ZVs�*���ү��6'��խ��D �v��X:A~���-u��p��� �)�`���K,���>��WwL�z7˜g.���?�� y�;�DM;=��5���Z�𭩽,�Ǌ(6�)bO�ج^����b΃Qڳc�/���l.ʫ�9��:��4bN官��t\�&�Y�>kH_��6	9�N>^�4�8��N�"�*�~R�׍s��Q�����4����u��Z�~�N��8�d:��ql��א\���<�ܶ��~�k����wq
�>��MLL���Z
z�������f�#���E�VO����4�؄���C��p�n+��f� DSd����}��!ӵ���M��?G��#�^:�f�~�����@Z�m�O4�Y�����yO�r0)E0���ʏ����V��(y�a�$���L/T����tY�V���L��c`@|�"X!�� -�W��J�[��MH�!�"$䚠�Sg��^�ۘ$s���w�Z�Fx�'��,�e.��:9����n'<d��@w�gg��Y���t��seK�aX��Y��Y�p� �|�Ε-�n�!�`}���S?W��˺Y<���e�7�(B,b���eu�l�z&(°�I�n�5x��S���i��$ǀ.���rbT��QI�x�^ꝎI����"�"��x�,���Q���/�K��ro�U!��:F������N!/c4=����rw���
f���Kwv�K����q$ߤ��r��΀��(�+&�2(�s�M��J-��-`"A��!���)�?Uڮ�X,.@|�D�
��P@�1�u�k�YI((Cu�!���}�
Ϛ5[s���M�Ӽ� ���]?KeH�L��N
��Y��QXilO�3��Ԟc_҇�|G(�J
������fA�xȕ1u��I��]V�L�K�_��@CV(swĢ�4�%���Q	�EHe��4�3����z�Gc��C��^Eb�
GS���Zפ8��?ׄ����qv��R@-oUQ4��B�[��h��y�q-�D�����j���#t��
e�/͒;e���H聧*�|PTG*�����M��ȏ㣴�~`����vɝ���0DڹBi�o����Ш:EA��5g��)���|�T{��TW�	��� �Z�%��O0���X��h�����6�r̩�V��b��n�y
�y��/ x��76�n��;{#��#�Z�V�ң�;���^���_<?4������2N��Į�g������	�9q+� '[�8��q��g����M
Pr'��]턀q���߭��{�a�"��N����.�g�;|���9�|��~/�[�q���&#bH���A��&�i���rkڱ�׈�uwn4IH�]������`�J��h+K�
���C�����}?�;% 2wul��Y�c)��_�@��48��8�ҪΠ")  %����a��������II=��wx��Cy��A6���R�����>���v�I�E�IȬȂ�I�;ܭ��L<�����V�	�,qc�!T�U,@؈b/ �+=	?p;�֥�#������fR�4�������������1�������6�Zs�&3C_o
U
f�j� #��6�g#���K&��' ����?�*?�\w����|�����_�S}D��#m ��T�~
s��D�In��X�>eA�
�����c�˥oq��[� V9F�\X���D`l�kgC��<�y�Jzp����-�-�����o݈�;�N�p볤�,�>g��AdqKe���\�N������������"�f�>w��ߏ����wsp+yNvO[q����uMR*�҃}�a�P㍅���)Y�b��.�Nx�~H��Z�������4���JmK�S���,�<�� iOkF���������~�H��?�I���5��d�[}�6 ��VuΆ��E%M=67��e�\�M��|QR�y%��Vp��$���L��,����e@4�4��`h�ʥ�P�\��lM��43�gC|kޯ
ı��'C�-E.5t4C*W���g��+��������kR�G]	�N\M㜀ف�,��%L��{���"�'oo�a��WRNWç ��� 
�\�E�u���2_5EM#>q��"��X��@^����C]@o�Up��D〺�5��/�w%f�֎�z�|���h���������`1�-���(3��e����!��V�\Z�P��s���C��Y�h�T	���Պ���L�e��JpY�i١nAj����b��L���<�<0r[����:,v>�'�z���������C%����͔�����V�w������=���T��<���`cf�wc�#o��M��+�LQ�=�~*fJ��v���$��72���6�����J$d�>�rc%�$]��4E�3���>6D��x;��=$R�ŝ������q*����^]������=�F�&��t�v��ά�閡�)�lov�`�!!?9.�9���^�[��3���c���_yfX1���V�o<;��O�L{�9�(�G�I��]������7.gbRʒ�{��"�@�g��G"���B`Y�j�5����(�	�ފ������y�~w0�]u蠼���B[�̱Csю���	��n�}3�m&B�z��Ot����GΕK�!�	n�S�����h��Z�����f�X��c�����aD���[���>��/��1�V�; E{~���`��bP8�.��D�{hDQ��G*��K�Anєv�j10P߇�6f�սb�Jq�SZML��`nt9c4A�]"�[�1hlr�Ж�s�ǫu�r��+�ʃ��G���Z����V�<���̥�*��b�q���U��*���Z�0k󗹎�Cw�/��'����j�E���F?��%�(SA�r#5&�7d�_`f�	�)��n1�0o&i�pJ-�)HR���� $\v	Q
!õZ��CQi��@pJ�N���`��W���K �)L����=�ŃT>����s�\?hg�rI�.�d��v�kV2��
B&K	�D�h�}�8��宿�t�:+����%���E�{z�7õ/+mb̀�!�M�����#���0�/
/��ޒ�x�x8 M;�2�B�����@I��0��|�����5�:�TP�]�����U�i#�ꔕ��5Xr�T^�
��k�P+g|��L��m�jB�t���D���R�ȥ��NmX|]���0Y``��?|�ܯ#үA�\.�+�7&��V��E1�
�
��τfIk'L�nI��G���Rdn5#�bh�aM�F����ӭ��j�"�(�\�w�M�3`Bޛ������b)F&;9�n���N�����Ałjع�S���\@j���F]����X=|i�w���e?�4mֶ���;{��O�Ǹ�=c>z�t
���%Z/s߲£9U��;��������ph��t��D<c���{1����a_:�Ћ���|��,�ɕ��2y���C͛�A�.�f �y6����oU�>����O�{`��=�N"S�_r���U� |�hT�3#� P����������a��$�8�ȓK{��'����;�7���|�R�n�4A�inbmda��*"�G�;	��S�hL�T{�	ȝ-.>Cj"�F�o��T�R�(yis�3�vJ�U�LAg�<���[
ݐ�t��	T����N�x��ǋu�{��_0V�K�[�|���1;H��$x�.���i��#L:�6'+{+��ܯ��%@�u��{��_nq�O�$�-�(�w�+�G^�T�����R���UJ����ť��f����o�x�f�N�賍\�!�3v�!��.���&�f�Q�J����G'y��uÖ�e��d/:����k�a�BՃ�3�軾��3�.��7�Qj"̙��e�����VÜ��L��dnϿ�q���UL��d��~ޣY�-��#��.y����z�r����\�^�b��ރԂNZ�(~KpO��L-B��h
o/�D��F%V_O��^,����!�v��Y�ZT��.i��a��E
��jR�O-,M-9��׾��^P��B���E�*�~ݛ�.%<֝��)��)m�d�|)���X��	�yU�0h }�����Ne��!�URQ���j��j�+�4� w%��<b`[�B���.�4�h'n�A�K��,���>8�t��:�V��@�44#�B��z�Ն_�OΧv��$�	��(+¦>#"/��	M�eO+$��;%�#��S��Q1zy��X��c�H����=v���1�	ӵ�z�K�����;�k�R��Q�^�$̀.�aȽ�m��rG�p�ؕ^� d�9+�m}T�_i�9�*��bW�o�Lr
Z�DZ�'���)�3n�D��Y| �_i
��Ƃ����U�u]�/Q[�Nw�K����k��P�Q%>�/%��H5�$^z�V��&�0�a^u�Z�<:Եg��|xx)8�� NS �f��
��I�X��N��((��fm3A0˶o��+��b�@�OA��o�/���t�t�vˣ�l'�Q����d������=8 �	_Z��~,�D�ڣ/�T�n�.��
%W�VT�����K�/��`��x��+�`&C�$kP�-T��p�����x�ǙI�y5��F��ڏ��o5 ��
f�ʝĚ�Cr�h��$��;��"T�V������D�J��1wg:�dۛ�vu±_�i2�,����b�F�)7y=���l�?�̩h�I�!g���=�r�j���*�j�-��ad}M�Iy�b�τ�n�����W�Jn� ܠ���0�õ���4M���T�C�A����P=Ҭ��j�~�G?�GV��Im���9#_��( 4�����x鶨�PgXil����9�C5S��
��C����@`J�+� �P���W�ay4�t�-~2����.�A,a�|.�!wp��jݾ��NT��M�f1:�x*c�u�|M�*���(r���©�#�ã��5���m+a��r��QAv�ԕi��x�5YG6n��_��{�('�)@�jZ����5�n�j�<iE��H-�P�o?=qu��7%vj��J�"GfB�������ƈ�?�b�7QÃ��B�u	op�W��ؐ��<��a�rL:�.E�Nw��n�Z/Wq>V�W���1�}=��{����N&�����Jg�Љ(��|�E���~vZ�'��^R@-z\ ��Q��<L�@���Hq�!"�~;ay(\����x���`�����D��� �;Mz�,�@�Ĵ�	��cB��
�ә'4H�_���'ٖtQ4O�o���T���~e.(�/=2qIw ��zd����C6{a"4B�Cb9p�(x�a[I�4��М[�$�}&�[�7��~��.Vq��/������HH�9�H���q6P3OB+5�d�/��@��>��b1ڲy�b�ږ';7kj�� �+R�̳��a}z<O���G�$!UM�I�Ƙ�&U$�	f ���m�����ܘK2XV��^bα5���r1�vf����y4�V٧���A�H��B�8.K@o�j�#`y�ٜ��5#�z�����x���Y��=#�E�~^A`Cj��^1M��������z8�3����l��Q�����͖X�)�|��O����I1-��(�n�h���F��g�R����Ϡ����;�<�bF��-�Q���_ՁHI1���)E[���4'Y���t�һ�y��J�(�Hb����OSA,:[��Hj�UǎH���Vz�&�����S��Iv��C;�r�������뛍[9Y/c�&��3���0�� ��Q�S茟x�N�y��)&W>��S��.�"�vGt�{lm5��:T�P?�#���UO�k�8�����j9��'Uc9� a�&�\Y4c曀�dv׹�S��g�E�"_R&�|B��j�ר�p2��u�S{�Ɵ���
!1�I[W��%u4/V�I���6EQ��k%������bu�ڹ�?E�jUvџ�����Y/�z�<���x�bL(Z��!e��R�p�+�b�sO@�*kt����ƙl��R7��������'�����7�O��c��3n(,p!�}��׃1�r��6�Rex�(e[2�Nߏ̺��d�3G=�f�v�(m&2���T���O�L34�@�a~.21��8�	"�+t>��_�����y?�`l�/��#�0�nf��v�(tZ���.s!��	ǔ���S�1pB�m�_׭�$�r�}2m._��q<r;�m��87�9�|~�bgl�Va!����z��8}����k*�|�{�1�kha�<(��|��=~R[Cu�a��r[��`>x�}�U����X|�E���]ւӨǇg|e"c
@
\v�J��D�;��bc�C~n�J�=�4���b�YO5�փ7�@1��ΔI�r�!R�l4���C}��f*g z��z�|.�$v�\���|y��䣓� g~
-ʜ�nݦ
�̓���
�0,�1{?�+�#���6D�\JU��B�t	�x�<��V�����,���Iث[�ep�"�G�7�V�߿,|��}�N������G�gݒw�[��^�h��I�-VY�SKI����y��:I��8o��,-��Ԇ�Т�!�t���ۢ^��=jt"68��o��Zb��]�[�����43���ջ�e��lGye8�:��a��dUۗQ(s�R��v�c��g�t��&����S<)����ޙ^�*�N>�2>��'��P�C_#���H�LF,�p)��h��Om$<�9�eY�Q/kgT��ߢz3Ily�ޫ�nBYǔ*�Xx�ohYL��>����z��V��5:�>ԺG1C�����s��졝�$8���bM���-��S�� ����85�����v>h�E2�7�\�ŧ~�"ZJ�3L�uj{*+�,��Ydr��h���ɚ�WI?P�L�ʫ�si�S~��Y6R�S�̂�N_�l�S�iuJ灳�`N����K�~q!$;�1�\�Ϛ[}1�,I�4�S[��،�@�l����DG�`�Hƀ"ߩb)|�+� ���?Sп�w�ą����\�c�Aνb�c�������ڤ��'���v�����+D%H�u�C�(���EP�~��1gu>���8%��nֿ<%��m6v��R�6bʰ޿�X��m��(5�IW�V<�.o0���.�bid��qn!
���D���5*�;^}���4N{��,�����?$*�1�J�Kq�rP�|���� ��j�ͣ�Ə��9-�B�3[jm|��^aA��߆�Ao��:]ú��;ko���6�eţ,͗Xcz�c�ȭY
��'��իqW�~����QBASJ�� :j�Z6E���)�EvGvR��U��&�6?�@���e^��:���	[w��|V-��|��|��t�uU�,��|�Z]��W�7q����)�a����;���I1#Һ�.�謹�z �����8��}uȂ�4au��%?B�0a�/J��<��-TJ�E���h�����)�W=sc��܊Vq�Xt��c�Rr���ݻtm`]��
G����y�H�b��?LK�\��vA#3��T\�i�f�{|/�i�=��6X+p��3�J�Î��]*�Sސn��@��og$3�qx[�h!�%#	�x���s��b���{�OJ�;<���c�M�R�#���Y����� �C��dE�C�����$|����b>)�#���o3�͈ӹ��jA�ɪv��.��9��@~��12j�c�y�C;B�A�L�
hx"h'��M���2d	q�Tx����>��ִ��4�$�]��M6�_zaQ�]���C���&�=��UI.��,T�i���Gi?��ଋaPwM�_C�b�D�8\�#~��E����D�8�n�|z����wv�$�!y��5[ ad��}3~8XE�5y O�^�=6�5�h$��z�d��ǟ���lH+]�Z`�����d	b�hn�5v�"2L���<�T|
�1�R�p)�%^���N���WI5��`k�?��Ū#�_F ܶ��F�OK�+��H��]�w��ra��S4�]�/Tq���T[�6o��G��"F�H}Ә��N�U�p+��Ō#V�e� 2�
�.JW���Q�V�P<e�����7wr*���>A�����R;��;��a�Of�T�,�_b�<�G�P8�9��7
���||�I����$ƪ?�8���Y9����{r�B��f�� ��1_C'f������]P�SG4�b9��V��?0)r�u�Icv���w&~�b\�B����%`Pv1 �ɮ� td7R�0�2��H�HXR������J��_2Վ�bt�o�_�Er�ظK���q�[a5v�da!A<;��5�QUx�M��e~�7*��q��x0d�Hɗr.��?mi�dY
�DYm�6;w��[Bղ)b|��7��T��%�#��v���ِ�T�g�@�]"
Wq�øg�#��G \��-$���!�dFV�i�Vbr�=�J�ծ��h?��T{�dE�x�,���s�U�>�0ɉa�Y��DC���M3mD�8��'0��#��I��3U�/&�0�<�r��A|���8݊q_�ﲈYW��˥N`r���[ �3G>�#+RxiLW���@��Q �w��!�A���� ��[����H��_mgT�4LMz�<�=^��.��5j@�"1� ����7���|j��?G6
 ����ʵ���gܾQ��d�`䲖RP%��%�jmz=�e%��XN,���Q��L�cRo�5��KD=����)V��!�r�9�|��y��+���~��1�����Z!1Vsf.���0mU�ϒ`�.O����a�w�}�S>��MZ�u6L�	0>}T*A�B�^j��Sh�TN���74��L�.�� i���w�ӧ�3\d�ɔ�̒��o�`���+�h�1V����J��q�7��]�k�.��^�=O߫�Z.x�F�B�)������G���[q,]q�аk',?)�@��酵�xW��t3ɜ�5K-%0�e@/4F�J �>���Q�7�e���v����Gt.�M�sl7�������bzQ˞G�6�7�m5oI(�b/W)ۀK/*Y�#x�f�������<wW�F���\^�D����.��?��
Ī��iq+��n��y`�2�H�!+�R;6��h�k�
�W��@|:�2�y��`p9d������4���I��''
1{��H�lS�֫��(s9��̠�Q�nù��6�����㡂1�QD#i�~�!=�짃f_���O��̰4�ǲ[s��:�x�f�[�\<�����6l��6���)�����A�q�%G~m.�
v��K�/�_��Eֱ��k!Ĥ�@����	1�@%F�T�SZ!<~�9���]H�k� �`*�7U���H����ۄuȑ~�r�l�]�g�v����"���M� `�Eėr[�;P��~�E��P��d6��g@4x�xR���+����+˺-$����G���E�B"'m�"����`G��yV���a��x +�B��u�#������:�h�K~���q�F�Ǜ�8mq�
.:]g���y��iS�.darR�:kARyxMs���o΍,���΁�NSr��ly�Պ���"���j�b��+o�3-�v\�hb���G8�O7��}H��+�7T�Ͻ���>�O��In�2T ��wG]͈�2�C��g�|��m��[��E����o����ai���B��7C��Ŕ=I�e�r��Eu{�Y�I����\Y������]��&6�����Dƽ�� C���<����"K|[�#1�a�ݧF�>5x�5#�os�~��M��'葅u%t��n������~���U����p:�B褑1k#ӕD8�y�üyk3���	���(SZ���R;P2h��ߟ�m�/�<���}��	�#�^�Nԯ#I���!��M���OZI��+wU���<�����p���ѐ�UD��Ͼ/��2?N"s��<��cCC�Ń���*i��h��y�h���5����Ru�%�@VaT�B���;���z�Se���Ec���^jK�|5���p��nD下{wK�$����4��m7D�p��E��{��1m�PT��|���ݣ��0�e��a��=���ڠ������I=�K��x$0P}h;��w1dQ����U�d��zI�<�fY�Ldl�3�f,��hG?��U>��O�f��
ma[��I8y|Su2?��%"ε��c�MӬ�Z;�H�U2�b��� ٱ3�r�
�UR�/=��8/(��׼s��45-\�̝�`�X���cIEHAXj�̸�F;k��s׉��q�+��_���fY�'�ʷ\@�I&�mdXZ�ksr���H�fv��:�36�X��4E"��ٓ�q�h����q�'ѫ��CWϒRZ�G�CcTNP����)�_捾!J��&a BZ�x���j��:H�����A	��s�����_nV����,	0�47�ǠoJ����G��	6��A�=�5��{�@�-�{��#���*M�.�hѪ�ATn%�G��'�aH�����vg*$ ���I��ɴ��Y�E�S$;>�{�Z�y[�6|����1!uQ/�G�aW�8�IR;s$��&I05� �.�����LTUL/����������4��6X�4��䏊j1�D}R�6ñC R*�P���4�[{|3��E��w�<�=zȂ\ߝX��Z��O�1�ln����l_O�4�\�xc����(�R��@t�@0iN�7�c21I��5d����d�pzM1�_�R�6��� �y1�O��Y������(�W�5��;�s�Dy3D�!�	�;_��Lq���Л5���#�"��9��q	�`m���C>�������F}z��>�:��dzP�q�|�k;����V�b�[R�/�ߒ���B�]�W�k+�Í����xq��������4ǭB��Ɂ����7�^[��U'R��� .�P��m~P�Ro��\�5�σq��$('ж٣���Ө�ʃ׸d�����F�w�V�H�䎣V� ��j�l�\,�`	��j-@��Ts��2[���;��F��A��~揆KÈ6p�!��N�3
�>��� �08-.�G��>��^�4��Y�L��qk�j�|�ĩ0;i:�(�p��+Ŗ�r�����t�$/q�I�.�D�LM��4�Z,��LO��r����i���<��1�j7�ue>h&T��i��
{��ux���?�r��(�ٵ)}��9��!���6��H]6yW��Uk�����n����Q�O,)ΥD����LD����{�7�E=��׭ )<�K��*��vG�k�ꬬ|�����^
s/��U-�RH�Si(����qk�"$V��V�a�OG�s-K�h�@�V� =7�% �Ր��V%X��%�|�#|�ҷ�6�=���,�H!J��t�|���]������I.E2��ڷ�D�0�(��ͭ?��~��n�(������ݡ+��=�h�d~D�/+(�{�)��9~z�_�:�;�e1��0�@���Uc0$�9&�
ګ�]D��_fil���0�1[r�����8���lY�Dl{���􍙘�~�]�1l�j;�L�6���4)h��H��-�l˼V�b'�'����.���B������M-�"V�s�A&���_���Đk�droC��c	���vҶ��y��0�M${�����t������TwK�!%�L�(��)�X�v��[ҋݟ)5#�%xƽ0{M]��b�g�3�s���Qe���y�a�w��Q�=8�D�X���d����;��"���^�0�m8B"L�uT�������xnQM���OOw�z�M�@���}�����$G�
���� �ɡ�?�* <�w��GbA����<r˴s/�`g��\1�&�Y�Ӱ�9��G�}��VU��[�����r�Ձ�w��0ے���!"��bU����q;>nb�g̬hx�q=�_�H�}���L⭋���B9?����8�ZN���ƒ��f�����"[��M�U���ӿ��	��/|�~MPNZV)��~���<�zWv�����8��u��M /f�3<3'M��y�_ô�.4�h"���!Y�F[��&9m_ݜ�#n!��O`��R�h�Iū����u��y����0H8jt�S���;ZP�g�c`��	�w�x�R�����@��tj�ZJ2�W�����ba7L���v��.y�.!��1*h��(�=~s���eK��C�L}��W`���YY�>�Ӗ_���!��djC��w:��^�V՛��M�p!��$|S�K0z�����X�ǒY�h��(��c#��Ou�+b`�n��idᯠ-=f
�J1�6�$��5 �F^[�4��e�/=����*�W���fgN�e���aP�I3���*��*��FD)Za����C�p��%I�0@
u��}�c�oh�m^<�o�[	����r�2,�8��}Ld��w�E܄j��_$�NW���M�L�H+�$�Kx��^\gI�iɎ��H��~��kV�Z'���TF<s�g�;�O�q��a"�(��U+�cE�{�{�gDk�/��}�8�䂸����L��L�� Φ��?�҂x5_�q{=�I�E��=B�6;�] _�b�"n�,Č)�pC�bdh��ȭЯ'h�	�G��	Q�������1B��9i�U�3��¾�i ��E�
������@:��+��9eX�Ǽ��p�= ��1��q��?d�`t@+��Лˆ���:�4���F���ßQϳ9f���!/}|�%m�3(��#)���Tą��	a}���>�Kb����;}s�=(�A!��+�m��՟簇�M��_�ct*2j���+on�#O9-6�R����c�̧�JpBy�{��>d�6<�Ȗ}gPn�dm9F�A�sh{��#%�ڥj��'q�e��l����3��~���l�
%Rg{�sbe;�����`�����c	����I�a�����1K�(�W�)39ͰX\�:'�=4�� �"�]�i!q6�F����� 4J��z�qgF����J��P.�%�-JC����{M5����_[�=�7^\��!!�(QP�AX��UIؤ�\ᇝ>S�60�!��K������1�-�O�ۀ-$���3�)6_�2I�����귲M�E�w\�wBkFh+L�)}o�UQ(�."n�>;���?��=�O��P�W���tm��dw�E���@���'/��ԍ'����#Cͩ:m��ӂx����/��" ����𓼥`��-�w��/�R�:��C񼼊���P�Ь$�N��9�C�H�q�L$��������u��v�R7�i�o�{\��$�����B%	��&J�D�Q85,&��3G��%ʷ���m$։�����k��N,.�}e���ȩ����dd5	������+���)���I���HHJ6�4gX97Xn*2�d���C���P�� 0	�T�1>w~`�xI���Z�F<]Uc�i��].(d� c���b}��Q���HǪ�)�t��/3Fj�%'���Z��p-�m*F<�7=X(.'�,`�1���nw�Ǩ�J�7�(�'�V��y�>��d��:գ�^i1��g�lҔ(�+�֟m��{}��h����B��K������/��ZM�eQ�r���r�[T��9g� �����n!]]?���\�y;A�p�|��-�lB����ZT�j.���S�pj���mա[���3~cf�D��g�#oȄ�\�H^�ɐN��@�E�c�N	Awd�(�����=&؏�;�$��PEO�2���쒮C�7���[7�"�����6�i�`c���캊N'�&���?����������\u�����ٺ�vSzF�>��� s�63L87z���Fe<�A:%�9v�3sX݆�6�gO�T���'ޫ��b@��6N��ᚔa��U��n��mO��#��AB&���{�w���	�=r�U�_�z���<mi�S`/�;�۱� <`k���]G�m0���i��g+��H����>u�&���v̔�Ǚ""��O�s{o�H�@�����0P��!�IgwM�e|���t����9 �S9��F�
*$�h8�R���hl�ja�3g�by���5�3�.Ih���'z�ñ ��@/���Q`v�6����X>
w��I�҉��pO�|O��#8��T��� �<�=у�K���E �q�}<:�|r�#�?�g������g��W21����N�UI��Q�嗳މC,)��>�G�ii�y���VG8��	���܄���P�"��A*�ǓzF\�d�6h���f�̵'A ��Y�Kq�C}e���%K(�`�wq���^I���1��~e�^�U��f?�S���m� m������j  ��"��Y�Z�8E�C�b7&����G ��~���S����=o�[�H�| ���q��k<u�w��%/~���6���$}ˀ�\U,�FE�/�d]�m�KHjg��P��ѽ�'����8�Bt����h�'A2kC{�zz�Jz��&ܭ;V�����1	0aU��ȗ��cb�u��K�>Ͽ���p�M��,|��rw��9��{����+[�/x+ů��bi,7c�4���k�Ǉ�s�k7g~�]�,u��Ѹfr!v6�,��ٴT�����{V�����I�O��[��u����N�oo�������kW�����D���t�����,�<�8yꧺ�=��S2O�ݼxi�5�v����\PX�k�+6�D��~��:�W �M<S�#t.&��"(�|���c�F�[@�e��}g�fDF,-�.������t�C��A0�a����x3���r;)��?56�����5�j��:T���\��m�Շ��=�l��l���|����ME�N�8���7���cM/�Br��ϏౖbERO�n��Z�\����?8����HK˧*�{^��i�r�՚�.�;�w(�/�S�	,��
(�RD��@��3���1��)�_}X���S/Q"#���<�uP�9
�!�U~�x||�C�o����<<gӝ�jo����Qv
.�^^&���E>����0�f&��S.�D3�!SE�n����D>�]�[��f.(�ѕK�0�ٵ��?/:@B!\� 5!M��>[/�X��r�;s,�4�$����+jݟ?��"4��,�qa��x��!�B��E�p�Fz,޼x�a��} �N�cˤ�ڧ~�E[1�"�R��?N���0w?�&ȺZ��VT��2D�e��E�� �˼�m���\Vf->�>��'5T�t��*��UӲ���Y\a>HNU#��JGMA��rm�CIz�|W�b�R�!=J�C����hT�n��7�t ��ìп��	�9����H�K��D���\�^���/�Ȩ��TpbTj� �F��?�ݍM�v�
����g4-ْ�ix����U���Ȭ�M$o*~erC�KI<�&�.� Du���X�w��a��?���7����6 �9.IƸ���/��w=#���@�*�Qʮn����9uS���#�����)^���w�Xf�yf��<�Uۤ=+���ւ��f0ޗ���٤��C$C�V���� 6 2%� /p������H�z]��󡴰������C��6�����:�D���8-�x�Ϥ�ۼg��J?�ew����K����<n݈e���~�, �L�����?��+B}���b�kl���o#���錿 � �@L_�%��`�W�>��#�ae���5;�%P^ɽy��A&g��}� �8�a�`��m�K���@6���g��=�' ��ˢ��֧��e�W[��.�@�Y/��;��;��%�����>��V��k�L�n���i,c�|�������
�R�N�S~̈́�����Y`3��Z����<�j^�#G�ٳk{�$p��o��MON[���"|Lw���dln�uuL~���&�� �0ړ
d���l��B��;�/㾂�,���@���WID5򏚸�~�O���mM.�!�������Un�Z�
��_���=Hǁ�3��_��Z �}Ac1���Ocxo]��u4jUңp_��5h�)"�% +�I$�G�#�����ـ�{&�����ն�Fc�����`�[;d8*2]���4m�'��A�62�_��t�Y�8pC�'��Z����9A�x!9&�������f{����"�=��C?L��ã�N��6xt��d���)T�S5� F�>�>�G8�0EM^������'Svi���f�[Aɟ&�Dʑ���) �y�ҧ|62�pG�G�� E$}�|����&;�̯2ʃ�q'm�sa��B�ۊͲ�်��:����A��?g�ś��?�� ��l:�͉݃g[,X�b��1c�I�|8�m8X�ڕ "��	�f\oR5'N~c1:{]��%��{�S����N䋱�b>1i�UBE�0�	Y�<��]m,옆�9���a���&�"�OE2;��(��ME���K�j�z�cR�G���no��M&�.�y�(�~K�ր��ܢ}՛�0�3׶ċ�`��*� e�w2zǺ ��G7���HY`�9浧(����R��󠜯��<���"oMm�D82��b�Vp� �m�[?au��
�!����uh�Zn"���(_�f��~�
WT�����+9�KPZ)�k@��IΞ�*��=�l�^���_2��9�UMr��8չqJ�j��)z��h���_*��惡����쌳���0a���7��'��g�{��*�H�IX��w�	��;X�o����৔d�zX���(����f�q��<~4 'R���6ur�d�!�PZz8pSfW���w��=�����L{%g>`�=�}���uL����A����ܲ�L��î4��J]��t��\�������SD�S2m�����-C���9����geluX7iB������|�d�(���겤�p����ݼ���tI�����ZH�p�\j.MK<=wJ_�{�(���������$�H�֔JO���1�]5���ED�8�?!n}m满	׆��ޑmV�q,S-�^��r�K�W!����1�[�"U��I�nB�y���]yG��%BR
Q����ى^K*����I�%�\�*��*��N+�y}��g��H�i܊���U��v6!`�]��v�!���!h�E�Y��F�0��k������q��8D��~�5��R>2��؀��N�ٿG<Ϩ�W0�J{0�� �=3[=M�֍J�'�m�Up�tB �O�|�;��{�_&h�T��qUDe��ڵR�/��3��{^�k�A��0�K���=qI�:r�J�O�/��9�F�2{[��-��� �&��M3#���@E��'\�	=Qk�J<�yu�V8U/�J�}@����U4��#�!���NKj*�T@?�cH�MqI}^I�� �����'��U�⾱�;����{&Ԇ��c�?�1�3Y\J��16�)�@A��Dw������B�جF�$�1�-��j�<�׀n�0�w�>�)m�vQ�<5��Σ��&A��j�T�ǫ�m���"U�V�L�Z;��ә�x�Y��,&��^�܎�1���r���5/�>�;k}���(�a�mk��b#��&}.�+;yl��(����k���U-�Dc�q�`$-k>��4����n�Ϩ�9�� �y����JzpW�ih;�����(˸��	�:���gM��������>3�Q?�P"�!!�����Sʝ����Wڨ?�9���洬3�3�eGnhv��D�x_O�:��}��
�`�*[8H���\��áK��pa{��F��e�偎���4�-��~H@����$��?M����Q㦊��u3��z��Y�_9�%�U	�PĈ�0�J���Qx��R�-�i������U��Y��=�K�0#����:��#�dŎea^�g�oD4Q��'��z.��#�j0��𯔰Z����K���oyx��<I�{R�(���~��?�:�D�x�<iֆ�.-�cl"�r̢�8�����ݕ�=太�p�n�����ysSF-h@�BS��O�D[�����BQ��Er��(p�jr���������oﾊ:��\��"Fj.?��cXd�k�1�����2ڮ����e��/�(�ҋ�omm�6��--ytX�l,�Gd��9�M&g*6�@�Ve>�k�3�]3�
D�]����y� 	�G7�8qa^���Ma��@����}()Z��b"ZА�n2�o4-,�'l���߮üa�Y�g��,��ga��T�WL��q��[���%Ϲ�SC+�e������ ��r=���Q����!C�Z��[�NԊA�gG5��u���]��C&@8��3�m��k��:�j�z5%���
;�r�'o��\f��A���PƲ��=�b�'��}����pb��S�B/�o�r���&��>T�=Eq��Ј�|�A��v鐂�7��G"� m�� ��S��¢9.������� ~�e�p/�}�};B;�H�t:��=-I1vx�t"��.L��ڻ��?	��ղ�>��1�'�S��g�/e����d#W-^��Ҩ��br��U���mQK����Z�p�k��Y�z���z���ZS����9�����I��j�ˢ��T��4i$	���*�3]����'B^�xd5/�У��A��&�V����N�����֒$�
��i|�ﻔ�2��hKS!�m�y�jS���Vc�K6n+�F
��*xv1hT�����l]�-EL�X:$�Qn�>8�?��W�ȟh*:��������y��ǟ������#q�z�i
)�tL���k:�����Lw��E���\!�Z Ş(A�V��$��m8��@�����U�0C2 ��q�[����vC��@V�S�ʋ�<� ��3���P=�V5��R��)㧨��B<m,f����>〿��:��7(�*��)���9f��^���7�P\��Lb(>�r�4Jۚ���iл�r�y�||���A6�&H�wp_�WF|x�6>>�9T�.�}Z��em�AI�-lC3�sK0S!E�T���	B���1�@h٬���&���.���^os	����]C��G�2��X�j�'��a)g�j:pАZ������)NV�/��/�f���dP�5��8��=����N�=փ����O���"�j������w�"���!24��Hbv�f]�j����8��o>�+�@$�H	��9�$3��)c���l�yK�����2��_����C+ph����4=�e�nT�4yz�"6]i��{���ʄN~5�xEqS��u�����3�����C��Ѫ�������YD�BO���`7�;��e$Ui���Z0��'�P�Ӧ"�s't��o_}�"�T�f-.#�=����/uBJ�H�̇!�.
�V��CX�H�؞=���{S��c9��&�}��\fF4��K���Ā���� ��P���M|
��pПL���3?ʝ�D'�l$��<����p�Í��R%���s�~&�,�+J!��O�h�;dd��y?;�ߎ���^��A��	n�=�U3��:���lsU��Kt����%��� ؒ���#�V*3����¸8D��cY���'�^|g�}��i��K��U_Z@M9bPJ��(�W�?��zߛ����
h�g'Q��U�+���.�F�#��#��������DB-�������8�����Ahv���},�'��l���Tb�Ы�B���vlߕ�@ّ(kW#��\�����ϧi���/��Y	!Dr}寓�P���By�_��6���5S�@�̛;�߉�ꘫv1F�c�ۉ=xE�v�X���*���pG������&�ϭI"��ǣ@�8]:�E��s�4G�Qegq�w_W����ub�Dܿ�4��p�oS��0�U�ά	ό?�{sġ�>������-�U���4���|"e�Bx;���:7tR)5�v��iޞ�b�B�(�"#����ͮ}�s�����J�Գƥ���@3�D�C7�S�n2+oHn��i${;G���,�j�?��W�st��hª_N�ǂ`{���n,���j߇OE?������zШ��ې|j4B�
|�>�M�-=����;ߍ0K߄-��F����ЯR:����acLi3v�Mo���I{c�i��&�#���#+�Ӻ��A�ٍ��<���y���3���L�'��FI|�kbR�nL|z$�����<�hx��x0!�/����;X�V��s@���I�)����Ck�-���I�%�9GGez�<@+�%��\�X4��0�� �u�^�ڦ�Bݯː���Q��kx�w�mc�hFVwd��6��#�&&U�	����.���;?2�a�$3X\݂i�J�!?l�A64�2���#�A�v�s�B[�J��Fأ��i1�88⟼BX�:[b
��2kZ�q`�������gw���)&`��H��>Jo��Yv���(����\����Fg?Q�hK��vG^�[��Ⱥ�BҲ���C� k��T]����X�`?�C3�(�?�?��F��a�������O��^�טp��|���[��.�=K<l���Q�TN� کj�� �BB
��.����I/��~i㧃_
�/�}��>��Up���8m8�\	&�r��	��i���aMc:���e��ЮM�R=%���PP�Ube�R���}:~��Xke�H���Ӻ�qbQ�hג�HK�����M�q�P���o/YU�Q�D4z���j�J:����n�­<�����fR�j6o!�Uh{����ݡ�Y]��e݉�|#��Y�����V�%_Kdf*�Q�џ�\�6D��:ZT�34�����J��G2U�\S'W��=�M��;�D\���lhp�y�n2�灃��,��;�lݯ)���@��
��D6ޭO>Q�W2y���fq*�UMΖiv�(�f�HU��!�����-�H�jYB_((b�����\�O�X��*JUQ�D��첨p��A�@��ځ�!��w^�K��_��-�렩�z}i~bc|���>��b�L��z��{QQ�T$�h�"�&��^���d�����bd���a�V7�s��U�8������p����Eё[@��ʪ��苛3Bmo.U��"J���`'<7�.��b S�n�O{םa[˛�z{��{�w8R�6���V�Uʷ���m`O��tq9�n��,ݞ��Tq֢L�a?l.*	a�� ��\;�Rc�[1��|���H��<�[H��jHsH�(�@��S9�2fȗ�7!��A��-�?�� Y4ӏ~t^<���������;>�a��-3�)���w�oz�uaK��W]��|�zٓ8>��_>�{�N�Y��쵐�Ptc�;	A!�f:;F��n�x���x���|�ćk��9�˩˿��<)�bTxQR�a�A_;�w�Kgu˕�®���m{�����r��>3�.Lk�l��S��w�,��`>#�#Zz���'������F3u���% ���$�DQ� ԭ2�F�`�@o	�$K�7�^��9�!b�t`���ԫVw�����D�����Q� �G,Fvo�*���x�A���N_���es���ps	��B�7��)ed��-��~���2��0z�1Q����b�(���Xv�	���gl3#kF���Wa���o���K�����I���iy*��-�/�Zh�U/�Bxh��!O�bp��V1ġ<��K">��G^�8'��|;?���e%G\k_Ӓ4_�q��f)#���'�HŮ��v��-d>�M�*J�zDR3���T�\�b A[6���0���-)	��6��Jօ�oU��/#v����R����<Q_}=�Bo�/i�]���-ǁ)tD��5��0�{��N}z��*�ٞ$�Z�ԬC����gKVr�;�tX�n�`�I�o(��������#��0�g����`b�!X��3_n$���*h<`Z��\_���I���SVWf�9�8ӿF'�����09��iiGhA��_���x�Z��)�wW/��]�a�k|��� !i�c�K��G�ꩽKM���N8He��:.*��ރ�R<B�_t�o'`]=?�4B�	�	��6X\�A�#~vp��a�J���G�?�U�t���]́�["Џx�K;�_�z�P��j�`��M���| %�!��c�IhHR���9��#l)º��������XS�5��_H����2UγMkC��s�{�]Tmv�:�����$��ixz�jFZ-����T�.�����:��m(g},mƘX�@��K���1^{���Q,���v������s�$x���}�0�up��n�}R��D^���^f�4��R �	~��#A7���m����9h_� ��0쥜����r��=����؂�e*-�:Z1l��1�^���f ��xY95�]�j�ؿ��pL�_���a�y���F���z~�J�D�{!�)9�r��Y��F�mt�v
���"i�BOD>���%_�G����]��{�|[�y�P���{8Ӿ��{�0��=;�Z$�(���v<B�?ؾ~7"!|��c�}_�f�j(]�.��g�~�*�U#��*�S�ŲR�GY�(<f��a�J@�i�f1��o\Y�*��EY�戄F7ְ��T���rb�M���/I3]���Rl���
j&�L�թ��]�:���;cW$�u�RkInF>�Q����m{��K\:�Wi�>dq�ǜf���?�I��@��`=��k��\���*Z�q
����K��hS�N���,��lˈh��� q�K�z���Tz�.	^0s��)�m���;�^�Ap�W�$���\�U
þ��TzN�/��2��&D8 `l�J�6�)XP(]�b�|O�ތ��U� ���╞i�u�����V?>��Xz(��>�2&���{G�wח�Hҧ�o#���}���^ �Ci�e)�ҟ���遜Ľ(�����VP?R�rn��^�����[Yq�Tm���������4��_q�8fi����w��fd��;���l�u���B�N�[�H�LG��X�0tL�^1�L�_A�ʁΎj�t���O'w�F�]1�"��E�d�󫌤J�o�.��:�	�p\7j���xFi�r�7����$�*Ϯ%b���A���$L���Q�â*�	�n6x���%Uv����Q�'���Yy�^���m؀���;��Z@P�j��J�΅�/���WX�������>�O����P
��vC˲)j!�6*B+pu�Z�ـI��q�l�̼n�=d��5��$S	��I�v]���!�lNc����?�d�)�����,�hy��M�}�sFF�j���~>�5'�-���Q��ܼf��:��:��G)|�$�������Dj&�\a�����Ln�P(LC-a)v�&6y
��w�ug+��0��k��6ݧ{�W���e��/���p"/#\!��c̝�;$l�eǹ8�x��4�`/���+�*���D� M�S�@�Aʁ����k���b�b������[�	Q��3Ts(�p�-qy������t�	����,4��W��e�?l�CM� �V")� S��^�vF�\��)հה.A�-�
�oq���d�aj�k�9<8����w���7Ax��V�	U�0$�i�5�#@�F"Ɵ9:"�8_U�� lᥲ!�f�k�!�2���ށ,2�i��ĳĕ��{|�e������k4��	�Lu�M�9��W��XD"N���X�Q�9!�
NE�*P��P����piC�i]2	"�#���AE<#Ι�ߓ��!3Ȑ۪����;��9��8��
47xUE;�U��\>e�����1�ĸ1�4x�[rm����G�L�J>g16��.cO�
���S��� Y��ҿ����H������w`�iҶ�s�Ba��譖z;��[B�(@�#��/,��c?/~�r�ۿd0|s�>I�mt��S'�㫦S2Xj��ߕE���ڶ���uzX�E�*�%!V�E���e�P��ʔUX�������3w&-�a��$�N������B4�����}%�	��2Q���MЭ�{*C���SW��o-�,O���:t&a����9ί�ڶ�TUy�o��4��[�k#���_��e����T��9��U��N���:��,����_���s��'*�%w����;�gȜu\�,&��GAu.�X9� ����!�H˦��V�v�=[D�/��i#��wJ��00�e��/a �ˀi�����ߥ���D�
��R%�(v���5��������w�h[���`�!�aۙ?{�:�*�b��yONp_��XPj�"N�<!�]���+.�7x��Y��{p���;p�vU1���x-$�<�L�a�B g}�[	���&��/��Gv��?kfe�;�Bc@�"f!O�Zw��XC��]�����<�Z�q�N�Ń4	��a5�L��@I͒��Wj���.u�O�xj=N����dyucw�IUGC
�wy�;OH;��P�/�7 V	7�#���WU��ځ�>tm���V]�-�g�b9:����
ss��ڴ���`��
k�V�-��[���{ ����1�7�d�t R���D�7�`�:Ӆ9�+q[��@�L�����20�Ch�&�*������ѽU;�A� ��O�f��ˑ�@�і��r����}��]b�+{=5<[�����5��	�u�D���"��Ff���g��]'fѷ� G.d��xƯ-1e�kgn"�$�۾�[��!�C�c�`�.�G�q-���e�!��g�t� �M2�{%){���"E�a���Yƀ�������>%��
mVA��z|v�f�'�#�{؃ɘv�[��?[����N���#��V�Sg}�M���6�?K]�Z�H_�
�$�a�6�޾:�43�A,%rѳ�������/�XU4��|�Dg�ߐ"*�7!t���]���OB8�A��?���(�m��M�d�##Hn�6=?'+�#:�77}!9��k��^��ckO�D9�>�w���F�A���a(���f��ͮE���q��V�M@�
=�o��H�:�h���3���b��DY���b��ԩա��0��?x����4��u׉g��{y��C��b|�	J32$g�R��ڤmn���N�瞓aO����K��e�	��o��p�e�p��Q��/�+�t��N���pm��5�F��|*��q��仴?���O�,�
�
����<I�W�W��s0ET7���{����%p��+�[<<dݸn��[��\7Ӂ�P��~n�}OcQ����ˣ��Uχ���-G�D���iC��,2���Z��'����7�6EI�;�l*#�K�*�^L��E��ԇl9hѲ�Э�=�#��>�RɩǸ=hj�c{��.�.{+���!U�v�K�՟�Y��L��ubaI0e�h�� �9C=�D'�z�-BP<X2�^�����U,J�G�z��yV�Dr�J�
�랅2�+�z���� �� ���{��E(��ʢ�d2��mY2��c��q_��{�p��rp�D)���Z.a����q�l���bF��juB���,*���ع"�Л#�ɟKӊ���l�j�q�cLE�HE�{�ܣ���&cv?�3���ؖ>m|���i�A ����ņʕ�|;�_���قIkk4�D����z�)�|s�[��~�*�zb�U�:k����6�u�]�ơ8��DJ�"2���oz_!@�*�<�L�33�$�Ů���;����
�l��/�p7�x�_��������m��OafX���>m%-��p?b	�D�����#�D
Jq�e��U:�SV��� !�ۃ���3��_&񛰱��H��t�ؙ��1K_�/'$*���G����
B���ˍd�Y�4�䲲��X+e*ރr1��G�xD�z�r/��Z����ʭ�-Ãh�L����̸�.��[PPڄ�C�R�HI1���Sd����?�1O]]��M�?����N���v�k")�.4t��(�"�*K��I�wAz�6�(� L���w��zxF�j�,�6�;���s�Y؃R«�`�X�-ǂd�S;P�pJ 8P�ڪ��)L��+����o:�q�S�  �H���8��fb9�ٱ2ԗ�g�Y�7�����M!�,#�ԝ���zh�<F$cY�¬�~!��������Shy�qg�ė�x�ӄF���C6��r��-�O�>�F�hF��H����k�ʾ��X����:y��>�cH�^���k�U+	|1�.�ڣ�`|b�+��ۏ�b�kc`b�_�m2��\���T+�i��;b�o��I�A𝨊����/N��
�v��	 Ax乳�ՐEQߛ�J7	��Sk��;����J��i���~�a>���F�xWX��`�݁��;��+ ����00�8W�p����U٬�\�����&Rnؾ���Z�R�g.NWW���]���m�������v������V\I-W�;B)@��֎��J�[vYˀсb�8���Y�ea�y%��,H�N�.��F�;��P�YQ��j$@��ݙ�$������>�Q�(��ul7���h����.b*ɹ�זzU�.��Wٓ	�c`ڑn;�'a�����9��3���#݄&���J�������i�X9�ّ��:�e�}�Zh��#�w��ny�N��Z`؁T55JI�
kG�I��5a:��P�������z<?=~��`�ه�g��Q�V���ɣI�`����+��̺ӑO�%��r;���x]Gv�E����8��|p���8�O� �A���I�d�Sx�9un	x�/<�s���r��]��2�exXm��M��k��v�.��)�m��r��71F�>x�|�?�T��Zic��%��+\{۔�T�ߎ	���4'�ޭx�b-�!�u���nM�,3�C�p;o�r29�L��Ւ� {��gO(4'�2��3��.BKvǕ@y�HSP�b\5k��r���Ӏ��Y��i+2�^�j���g!^��f�S!�X]k����\
f(i��c�N�&��R�oH\�ͨ0����3���Ƥ��ޡ���%�y/B��	h��P�q��*����BW�a��H�����^��Xu����!���*B�f�̡.���O!IV��e"d�~f��^;�OFU�*vzYc�"]+D�����1wo���7�E�dI�B ;�F4�K9	S\&y�^�U��fx��3�Z!���^I^�n��a$2T<�O'��(�k:Tm��<���2[CP�_� B=���F��΁�飌�r�Yv��ҁ�������fy��ۙ[ƣ�������=;�-�@9Μ����58=�눙�vqrx��J�t ,z�#��L��� P�+v��&�����4i>h�0n������'�8h�K&D��W��`%�Đ�բ��.Wq��m�;Ν��{&	�F���r�=Y���b2D��+:@܀�\F���V�'8vFv�&Pf� �l+��#�ڊ�{~9�mTh��b��ݱP����M�4�%�|�b8z!�F�ַ|�h_+0H{�f��x΢���]�^�_7fa���z�*N��x7��-ȑh�g��~r?��te2.��ap�?"�Mp��I �ꛀuJ�A}��W� _3Ò���\�΂���Kb�ˁ�L���5�r(E��`}&�xр�@����p.���r�)%��1���1	!��~ҡ?��c�{cʬ#�
�RQ�z��$ƫR���/u����22�����1s#����s����?�������OZB�z��Ј)��ث��6�(��Z�a:�y>!��:x���v&i���~��u�k~�꩙?�k��#@�f_q�%'�'\��P����/]��%�_	��?�3P�ZV���Wޜr��� 0Zx֬���O�_���S'CԙҰ+_��Q�y䵑;����i������tjӺ��8�1�9�Kʘ�J[�t|��2Ϛ��̖�ҝrr�c���{xV0������}���A��n	|�
��`�<0�'�^O�V����:���4�.6���p8��+�hƌ�z3�$��l��̫�u����6?� j4}����*�ϯ,�܅dw|\Rj1z����h�L��,���ȃ�g��"�����	w���q<S��{�4��eKTPt��U�"�2���2���?;�����E�鸳��R�Ж)M��5���؎/���ԑy�c��~[��K�۩C��i���D}�F/O��^K�i�CÀt� H�D.*�]2'Jd�mz�8�K������EjB�.��ݱ��f�`���vlm������,O��;_�+o��|��Xjh}*�c����%ê���_��{���v��j-�e�\JO0�J���Q�U�{�
|�?���T4�g������N:H�	M)���D���Z�wӆq܋��gu��"�����k��$�g�&^BI����&�+jf���"qy�I>�(}�m3�V��M�<���������חyh���L�iy�]9�����M�؉�;7��f�;�D�v�zh��<��%������䂧�M�M��ƣ[,�U7l������J��z�e�Uc"֛�������Ͽ�~�H�T��>E��8�!-<���Qj ��%t9���ڵ�*C�-��� ���B��*ʹg�1�;����?�񌬆}n�<�:�2ZB�Wc��#���-�Q;���UC���5�r�V����J��� L��=�:�8��LĐq~�Bȗ/9���_�ٿ���������΋+}@���'�^GF��s�L�6��9gIVx��� �����<~:&.2>a�Qz2k��>��\���u(ҡ��M1�&�X-�Qf9�I�p�@�̗�З�|��'���(�{��#��>�� %�hz�Ӊ�z��E���.��nQwbT� m�-�m��Ö�:x�1�@�GPK_%�����wFh�D�Kas
���R[����އ�ZwT�]Cj� ,q��.K|��-߄�9h�}hL:����9��u �z�ԤɪD���_�vqmUdם�ʞ�G��d�!��m׭]x@�"�D���V��5��+�W,�R��N�&�O&I���T�w�<G�]K^Lx�S�_�vy�_�<Kj#B,%�E�0�A!���?���G3������	�=A�̄��'W��dp�?�z���U� R$W��]���E0��ؿ�M�ZL��`	.��ÒK���QM�ޮs��읲2Z��%cJgz�$�.>T�P�=Ԯ4�y^�px����}��b�Z9���7& �:G'�VZ�:����ó�s5wA��n@��#qv�'�DL�<�������qɤ��r��2�i�)�A�+��@�Dx��ϻ��{�!�83��w`^|�ҌyB�1�j�1����Ř��ָT�{���Q#�U��S�a@18A߯.����Ұy>VP2��H@�c-.�0U�Nq��OE��77)ç��b0ش�a��`��wci�C�q�NOSG3����5!Qn�=	���4A��#}|�>�kY��q��9I@ZBHz^Q�f�o?��x��ƌj>��p|�UW�=��)�Z�;���x�6�L<�����ce�'�H���ov���ڛV�{k��W��f�qÙ�\~��J8X��z�_a{-Q����c�z�q�'��Ä�#�fW-iES�e���s����y���"��t�:w�F�9��|��#R���ĵ�bXH��0�iꨩ�`xS�i\����v�4K�f<��-�`P��\#��eŪ��=��q��綟���e'M%�(��28�/�C ߻������q��f�f�/�?r>Ҟ��|����.���*'���^����׻a��M���㡥)��	�կ�bq`G#�J9�_�C�����n�P�~�X9
��i��*cc���>��͞��G7a�V��E���kZШ\�ɁIz뒀7+��.��}2����Bk�<~�z#$��h3+�U�� ��N(	�Дs$g�C=vQu�������^�Ӡ�~R�V��i8"0G�s���y��L���\ǡ�C�c�0�Hfo��((Cj*�{��v��J�>������2`�]�!�F�F�Zv��j"�~��R1z�#bx� �7���Z����Vë]y�WlcY2�����S��$�c��6��%Ac��5��B���@��G�+�)܊?tS�%@�J�P�ֺ�D9�8���`��Y�t������� $�`����ўz�rY��	R|�LP�Il�7*����&�#�L�5��-��7K2���Az�h��}�#��ᖗ6�����:4 �omݺ#�	bs}��8�~���e[Pk���\��%S=_���m![��K�����t�d���LT5�&A{�t}T��>�r�faK�Υ{#��Dr���.ݹC3K'�p�5=��=2OE��D����<�]KFO��m�VQ�G�S��N��nyqv���;�׻��=]������S@�O��T�p�.�km�^��Z�]F�0>Ɍ�-����;�:I�cIo����Yj6h��鿜0/QR�p�Z�n!�+�vM/��m6|E&W	�4��WI��yq^���D�����MY����d*7}Esi݄٩J�]tT���*2mB���G11'��p�T3�ts�C�p��tT��P f��r�Paꃱ^��n�Q���8�bJ����ũ�;��*���)�opp������$S�x+��K��S�a��Sԫ4(�i����,���D��ɘ��	���|}Ybp���[ՙ���H� ̎�21E��_m��C�0����ŹqXw��ə!��GXrp�q0m!`Ta{ȓa���ɧp��l��"���c�8�2\�F9U�^�z|q�s ����!_��< =�U�A)�!��H������c)���*����71|Z�����r?{��
M����ܧ>|n�
]�,I�G渻��_޾�Js/B��g�h,�$I�[�t#�cF���ݷ��-�*=��O��S3/�1�+�c���)ɋ
E�9�S�(��y�����ɝ3����P>�J+-�߉'0V= ��*��/��Z�s��;��4/�>b���� ��xM�# |������i�C�9�ރ�[x�0�.k&+o���9�/���SD�Xv:�)%G�EG,��y��]�s�=yP	���̗�|
�ojM�W֓�pʟÎ{B��z������ M��;Ku%[-�/1�R�`a�9�:$d����V��~>��;%@pŧ� r�nQ�|i��3�*�8�$T��پk�GS]��������V[�%�v����i�Q����X�$�`��MO�5_f2	�X�&�@�T��ޓq�}�-V���n�hi�y�����7m���#4e.yf��[�7��}5%�V}��$��+Qe����U�<b��lWkQ����E��i��J��uG\�� z���h�{Ϸ3�}څ�K�0�*��. &�L� |����W�S����<fq�<�P[��I���K¹�X%	KpK˨�N7��,b@�U�'S����'�m����o[�S�}F��&�[�~�mA+d&�N�4�~Cu��۱��y�e뛽K��EqY� ���Fu����q% ��ʩ�Q��J�	A�{�|~���2��1���3Av��u�t��L������>���q8dw���)�ݲ��O"�7tT �r��t-�I�����y�l�K�N����}�^�MM�,�DZC�!^���j����$|�˄(����<+V���KЉ����K?j�'�I����3'��v!ƫ2A��ȻBSEH���k��]Ͽ`�\މNf+�Ԥ��P��iȩ{�.�u�!S�|�9����{sv�-x�Y��7\A���;��!]��!V��z�`��Q����������"�FȌ/�3���DF�P|���hJ��#�*a@�`MR���
�!��3(�*��YsK!`��3C{���B	E\�O�'�KUm�ޢ�$�M�TkN%q0^F�_�yl�`��M���S���yO�!-�<�+c��a���i���s���qj�	=M�37�~Tz �}M�[u�X�=��lަ�xG�0�m�ѵ�xxC���cR���F��Sjr�����L-���ܴݞ�niv�Ax�/s�aNi/��+�3��g���l����������s[p9'�*���b�	�(;����R��x���G�ё��`#Q���nM�5�Ôp|�^)hN�qg2ݻ��уm���M%C>���8w��\x"�k�
P5V����g�١q���	D��h����
\���s�~����}���s�S�����`�.=�3��G�o)-�#���6�H��Ñ�ٛ(���\��ݸr���4��K�� K5!�l ���A���F��.,u>t3���_��`��ZE�ܦi�r�	\�@��H���g�L.����ح�lP�;�3��VL�Y���!�x%C�`8W����+Vbj�IKpD	2co��v���H�ƫ/b���Ud��\�M*�ލ����#�8��0��!ǣ�q��@1������<���ٍ�`,���o���q�y��[3<Wn���!��V20��2pTn��@�k�W�;ea�7�y:��v�&-�FQ�A�E�a�R�pb���N��p#A��g�#^T�&��.N�ؘ`N*I��0e��?�LO��~�οNV��R<���Z��7^�ùz��@�sۘ8��X�L�b�B+�F�m��	�����nS;{E�I�.��M�p���~�þ�H2���X�}�|/#�ˀ�P�G���ξ`���$��z}������[Dû��g��8?�(�EU��s��u|��� �O���+�:���%�O���q�'�,l����	Ʌ��5�~o��Z����X��])��Z�\̢dOM�x�g;0���-�՚i�:��:��%!]��������g�j�ko�瘕�D����s����p}�'g���ġ� 1�FvD��<ULpz�w��.�LYJ`+��̲_�Op;�۝���s�=�O���D	'y������T�����wW����y���l�O�Jn�Ѥ�2ˀ[rf����g�B���>d��S��Oj���3E�I[�V�a��	�ސsi�?D����(��ľ킉�.�Qy���:vK<��P��3r��cb�2� �_o��wN�.7�o�p��דl�mpI�7 #BѴ�����ó��>Q��tO}�(׳V �w�}�C�n�� `V�[�{O�KÌ�qw.<����CG��^]Q:k>A���h����=:� ��.�`�H��#��r��&�Hn���A�K�F��G��U����UBS��@QM�Z)7l+ἸV��%{�Z�*D5�_S|�*Ұ_c��n�+�����dV�-�ZiY�ӽ�ٍS��yoJ�z���|�p���M��o�ܿ�K|����%mSa�Ҧ�WP�K��"�z�-TqUr��r�0�XF�o�����`������C>3z�qx��A�v����{}�u5�Yl������X���0AX�w�?2�B�>�4�[~�����>=!���WC�ٷ^�?�oљ�v�,��I�]K}������R�������(���yѕ/�I��������"��������8��5��K�j��a���Vƒ9i��aH��x��	�͚�š��;t���ױ��z�|O9۪��8�����GIq��\sLy�Wn���/��~�5�
����E�6g�����GWb��~6	L
��C�����)�P���;��0��.;2�:���Ꝓ�c�g�{iD�HtT��|@_�p+l~Ws�&?�:�#���=?M���5�Ou����>�?~qo���'s�THH�`���6.M�]�GG����Dnv��.�:QKU9k�bD�Anm�.u���W(�كfo�a���2	s�zJ� ���Yk��+�2�A��!z����b��c\}`��`�P^*��禶I|�曷�eWf������Ao ��{�ԥʼ�.v|ŋ%��ch�g${\>��(�h6{g|�|��9�X�F�����g��qv{��?Tc��`.�`&�_G�S��c/��Ll�����UN�m;��X�[��OS��'ӽ�>�n��mg 6]�}����X�,��W ����g�%_l�����jI{l1Ov@���Fn>tK-1�ta�Sb��Q<��pwU-���$�9��NfJ�����b8ȴ���g�ö$�}ٕG�@���v�-��f�o�%}��#mk%��}��>S�x]%�g�����F`��i��L�#X}�J�V����(ݽ-�>i����ۡ��'�<�� q�on͟��z�� g�C�0�7V�	��v�A�y��R�4�P;��J#!�?�)��={&�H�&CI��:�
�n�3]س����d���HA,�[���'oh�[�����Z`���	;4�2���[��gߚ�KvK�́��X`�I_$����_�$�d�VĘ`�ɵʶ�fh0��{�3�ã�\3Z$rw�]��Հ����������'��Mv��@,M�&P$��� Ma	�GX��N����P�>7(}�G�¶�"~oܐH�W;�k �΃A;��
��ȣݫ�/K]nv���c��U���bqc͌Z�Z��b��1��Uv3�gE�{o6�QKQލ|��KM7W�8�	qS�^�`ΖO�`m��Au�n��9�y���
V�(4s�
]��{��Vö�p9<�M��ۥ����#��r���w�.v虽�B�A��-��K��&���,c����$
���yY�V�~�1��%/}�;��)���ˤ^�L��f�h�ӿM�]��g͹%h�I2֘��:U��-'�h^�z��%5�-s^w{|S� �Xu*q� C�f�}�Y Bx��ةk��XN���.���+�c�:��&]����_k%���|��� +��A�d�Ή���(u�[|��oT�<�~���#��]��d)���1�����@�{RxPLiB�?k���J}'kO �g��@˓�*�Xa�*0�
�� 
7(�o���ǹ��`M7�M(���3�H��FP6l�8���ɲ�n ������LZ��3�]!1���GC$.Ò]��9x�7,��y��a%���3� +`O6�.B4V��K���,� ;�����n ����/���^���d\2E����(Yس�|B�Ж�
_.�v9Ĉ+,�*p�p�C�՘T��m5�4���8��tङ�  h!a��ʿ)c٘���@nK��.�Kgr;&tV�:C��|��J�p:����v+�N
ˎ�[R�[�����6^�4):��O͟T�:)�P2�Iq�`�,��%�+(D��R���ݳ�S&[�%�@y�M&0=U���B��B�7'|�1�l��a���ޭ[Y��e�Y�X�=R#\�'�;�����c�!���Y�,Mo�`�9���Bs��$J�|�)�ūD�$�9�H�$���WJ�Q$XN߮,P�M+�NM|X�RO�[y�R� ��t�b?Җ0f�� 9�8Ly��$�8�Z����Î�������ԿgfL����ز�+g�y�PMZ���.�]YlO�7
�
-Ȗe��3-�7pP�
�n�a������z������'Ԣ"\��-���ؗ#�E�.��oY����<k��<�==�Z&|ĵ���΀�wC�P�)'7�bfk�S� ��p2�,��u�PYh�����	~�2���4�6>�$C�D�=� �c�S8f�Ϻ?��li���rr��}��Mj��p�v�ƨ��q�9F97��Q`�D�Ȳӷ��wc�),����!�hI>��fk|�X��jX�$��I����?r�M������݇����8�����;���%�#Y����S~�ђX}: �S��N�M2���il�0>��0%���B�t��x�2)t�6��h��d�������I45@�<9�_~���.2<>) �=k�R�ZԷ����*�lzP�y��+��dӇ�9��65�y�t&��rY5�D|�?�,Ɏ�1q"�Н���̡������{D��[�k1(���!7��̠z������x3�W-:�"�n�Y=��;;%e��I��4�G{�;l��)3 �{��?��H��h�n��Q�D"
XB�s<�єq��-�(6��[#�T�@Gg�1r���u1�"K�=#���&�«���NZ����	� 8���RD��S�K{�MS>p���N��LC�NU�`��=���48�^}�7����8��L�c0~����m]�����ԫ��>�n`v�8���_0"��2��!�2x�G�Wp�����g�c�i��A�k�0M<S�zh0���jus�P[�
H��Z��K��'��XƱɛ��⩜j�9U5Q8��:��غ��K�<,P6�V��m������kRC��AS$��E͇?P���:��_�fA�-5q��_��蝚�Ugj��?�m2K���S���L,B�g�d�_3|�D��y��K�"(�c��s���>�9״Mƶo����3mE�h
7�4ǔ ��n���Q�I�i�j�b������l�WW��6���3P<E�Wu�p�f�o��ʬ��9���֌�1��#U��(=^�0{ʖC��
ʌ�O�~�O{ �� L��p���+K��;7���w�ޏ��}�3��x��#�	M���``��:�������KN����B��v@�U���NT���?g�BK�31��5����*`�ڜ�8��ɗ�C/
�:A��z ['��q�=>��-��e��������b-P��߶Nr>��qh�I�5�om���u���q�G-��Xm&aڕNY�Z����_��1<��X�n�b�����% h�u��N�x/o�0p@;{�h,n��ow�&��a�ȗ�A2,+a��B%yp~>�$�*�����]N ��`�0���284}���|�~'�np;���4�F)�3��\ �f��ɰ\����F����\�{�W<hO����"�9�Yd��^�9�T��'�mV70,���+�ʩ:W�CYrH[ÎR��gŗ�Z&�5O�j����e�\j[`������gګ9�)���uU#���4	VH�]��4]�aFm�I��aT0��N����� p����#������JvF5��= �n!��w��}%H*ʓ#�"�#I��NtN��(���V*u��ɝ^�e=!B�4
��o�8�D��q)::�l�f|S+ժf2ÿ�/�
UK_�A�Q<�k1w��9(��.�I��`Hx2�5��g��D78GR�n���t6�a;�����I!����W�56trZ��5�"�6��ri������ �,˻JSϫ��
O���{�}1;H=�7h-��)f�O�[�+ �N�ױ|c��<~����x\>Zʟ�7�����7]�-y�#�-�yZj��&�=�/r+�{&4C�3*}�^��+�Yp��NHp}��h�>���q\s�'��wU#��GϪ�$Kj��`�
�O���ݲ�w��u�,��D=̎nE�]BT��}
�4�{�4�S`���Pdj!d��	��S
bD�|���}��(�r�1aFE
�F��?�ѷ$GǴ�y�(�Y-��l:&�{�)��ix�z�6b��H;1��ɇpH���u53��ѐ�"^��&}��bx�+��
��	L��}��#2õغ�G�Y��hj�~�>�f�z@��,'UT��9NN�fs�k��Sq�ph%�%K���!�B��V�[������������o�O^S�ETnr�{vw T8����N^րa3~m���iJ�RM��ho�c�;�<�Ħ��o�������z�~8v�K&��K-�X���z}�2{&8� ��&��Jv��t�A�z��=<�N�tWR-��^�H�Տe�n�0ZCįYDF���m�&�L��͏�2$�e���y�ČH�#�-�^����~��g% e�h�%g!��up;�su;���=����-R�p��2�a1���(����"	=��{����̋����c}$�����u����˩�\5��2	CM�|�uJMdȏ��4�lY�@���g#�N،��Kd��?ӷ,1���9�t�4����p�j�	ij�w��?�HGa	��ңw�0���_�>d����҆�����N�2E��&�]HsB�b"���܇��;��Vh�ī�4ː]Z�/��Z�̽B��Y"]��� D�V*����=rDFA)+��Óm5IG~�6�$��
�yE�^-w|�}_����[�C,Y�0�$k�l��;��E�u�?K:o�Ɍd�!(��A!��|D5%�h�?;;Rx]诡:y��0��D�q�s��V%���C�z�le�J�,�=�8�7G2G��6/���P����{��uoC��ڬ���o4^�.�%.	{�.���Z`<Rl��rf�a���Q!�6,�� ��Ȭ���z�����$�@�(X[s�wG�"����L¹�Y�!@��Me�d|dJd4�9�����Z��o࢓��}Y�L}�.�����,dF�'���2���#kl����Q!z+��uT���mP$����T��@� t�~Y˓�x����KL
8�n9���!�]ʃ��b�#g�B�g/�hЄFB������W���ǸD�*�ewH0K\Hc:�A�E���E���3G~S��Wl�3尙��f%� �hO>���ln�u0ё0�1��n��:�S���U��-��lb�՛}<W�gn�I�&b숧�Xr����<H���{��ǳ�k���P�B��^ ��q �&�(-_	�5��<ɥ���P׊b���yJf4 [��\Q�tꮊ��P���u>��2d�=-�KY��P��uR��`-m�Ȉ�����m�Vxܬ�y���,,�k�rA�a�=��k��70�������i�������s"|�  �L�_�R4�[Os����(��_<�3���M(�(�P�G�>�h�?�j�M	����dJ��I���w���۰�V"�:�GX�6��>A�*��=Q&�N����b��PR]���}�p3��Q�י��) �T7������C��cK�����6�����-}�N��ĞV����pK����8,x��ҷ���@Uı8�A���L�;8�<�떠-l8oɪb��+S(��P����V��2��(M�R@g�7��t	���Ϳ��� �䷽��h$��{���ܡ|KB�4��X�+}B� �U$�$�y��!�B/��d>�0�|����*vi�	}Ke�a�*G�g��]�1��#qr��Ï*��}v�q�Ⅺƛe��#�hWT�M>n��Z$��j�7M�Z���6]?�j$�|�4ۡ��,����������o���M��
6�I��<8�U��?�E�>]GT߯V��?a]�����h��pY��?�8�'m��o�?�+R�����6¢�[$�9~�$MUdt����(�:>4�.X+�MR���j�a�[A�r�'���d�L�B��v�n̮�D��MW��
��ј`���&����t��R���E�,���Di�c���7�X('��e���r�w����2��&#��c'E��)?�UQHI��/Ƴ*;����l9���
-�=�
1�g�q�3�}�t�����".����%���-#�ط�^���*.*lq��2�������Lѯ�:�W'G��l���y��X����'f��]5���D��"�s_�r�'���0��f��$es��-�������ڿ�ID���]6��&�`� R�C�u;՝��I������G��֨��_�C[�=��f.��XAV�$�.� u�tA+���&G	���г�,�&I�S���[�F��*�̚j�eW��c����DZ��F<W�q�������P�����M���Mq=LR��N!�A[������ ���.q*rBm!��ܲ8�|8�Q �Ѡ��9`������ky0�-��5��`�.)NIڗ��uQ�٦uߝ��H��Yt��d�~�ȑ�����#�&L9q!K\�d�'�_r��Zwg���|^�a.�o�����z�/d�A���j��T@P��K.R��Zwi�6��Ȼv.�x�槅E�&F�����;Y�iH�ߚМ���R��C�a��\r%��â��j�-I~U�z�r�Gɲ����!��}�}i�b��e�T3�F5�j����>��Ӗ��"�.����ي�S�nMU�	h{�����*���mN�љ| f��y�C#L#͢3��b�j*�S;J��q�0]�HY����7Q��pL9����C��D��?
yם���� &S'�=C@�๚��7���� ����+�1�Ќ�U���&����2Ԍk�K���ݞ$�v��KD:eE	ݔmyH����)��,9�4���n�b��a��k���� �a�;����-b,��i����K��R�F��6���-�fN��H���W�t����e��ӳ+�� /��cQ��U�1��Z⍚��A��\�,�q-��
x��e��K�ჴ�Gd����c�7�G�P �n�����
��W ����)e=�6c��r��3�����C��;q%�k�mQ�%P=���vf�б����ϝ.ʾc��`ݻ56��o���Ba���*,�0�<0D�����y��j.�a;�&	��t
�,?um����d��_oe�=�J2��ռIQ��R�;��o��#�|y>�:���xb+��/��t�jUD<N~j,&���u/M$���@!sm��ο�N��\<�$��+p�҉�� �`�^�\F���v7��	�H�HS�[�o�Y��B]���/�n��K����N�E�`��-ձt9d�;�r�+�k�j6Y���îvkg�I�p�v7^�G*U�K�T$�I1�����NGR�\��f�E��Y�qڻ���(���Ђ4����%��O���vM�Wy�  & �����`Y���:��{����R�W�aA�+x�~V��_�!,*�*�
������Ba&dS�4��������PU�������Ҵ�Q������9T����j�����DL!�R{��'	��ʜ�q@�]�9@9X�G�Vލ��P;:·�U:\��i�y�:m��t��C�\�-&E�L�ìf#��&<[`9�u�����E��OI�444ͱ5C��,__G����M&+�D�Ѝ�T;~{��1�P-�Kx6&~8g$�
e��T�C^���.8���9����6���l$A!F��~-A_J�Y�Q�@���(Ŋ���
�,����$[���՞�R��wfo��|q{E�<��8�B�����W�%�I�5��݈���V;7�nP�藃]��$�v]��6c�C��p��8�J�O%�/\*�^Oǲi�lA���iv`�C�&kҪ���1��N�ڳ��S�)���=G��@p��տtH�m�$����q�sz�G��ǯ
��n�߰J���-ψ���q �Z���3S~�t���K&��	��������>�$���C��W3�Vӱ�.�^}$�S����x��M�ȿ�>��P.e�D�������^��m<?ׯ�k���1je=;�H��6�~Z�qz7d[��y���T�D�˶��l��I���q�z5�=ީ�3���re��T��J6۠�����e��5�Kz:����NPB�*q�Ä`���]uh���z������^ԝ�"ǭ���t���r��ҧ4�p�B��)�v�}eԴַ�e�y�`>�qkB�.�.�m��d�ĝ���)�ju���4���
KE���\�w�����O|������m�#���f>(�E1Q�m�?GI=��ތn�V�Q-�/ ��?�����+n5U,�F��l�+Az��6��4��jh\K�6I5˪����zM��d�<ֶ3.�ֳ�SW�]̹2��b=�%�~��
}/�>Z��)L	I�
�l���Y�����M $�	ed��=�z 8 �zք�����1���zi�g]5������4ǋ&z�	@r	��[e[U�/�{K<xβh���r��_{�CH��UC��Z~�qO2�R:�CLi��=M�8�B+��:��_�E�N]c���N�m�=���"�����P���e
_�S��Gr�W���8��$O��UR�����᧶ΟJ�܌�ԩU�����@q�M���4>�j:ʱ��2���n�>��N�^g*�
�ޠ|D��e�g��m��s�ȡ�8��k�tc��K����o�w�U��%��m����l5��ԅ�.��5���}D���<���lK����;qQRpTM$=�J\'d����tӥL�X�A�:TA{����8��c����_�,Ж���YԆ	l��Z�_Ŋ���TP�y]����<��|I������J�¼n�ԍ�iO�G����d���/[�AB�R<Ƕ$��s�WZ��~L;e����J,�%�Ώ���������U�#�����L1�E;��?�/�Ol�=�P�I̻W�s�H��[�b���1jZ��m��I5�i'̑q/	~iⳠ3�R��*��)��?W����󟢬�f��c������1��[�@������[���RK�\c�x�P ��H��c�1�\��Z��h��7��e��:;�"����=�OD�d����<�T��Q���&	�"�I��v�=��I���UJ ����<S�,�h������VΨ��
	J���f5vb�K�!�{�џ�R#e#C1vG��mʤ�)9W�M�����]�9(ژ��ٴ�S����@{\�Ś�vŢ���1�Z�^	u}��30�#ɛ=eZ!P�Bx��4K�J>���|�UVrR���άMK�f����dd�٘�U�C��l��]<;�7�)�c�B�uq�����5<�`4�Q�]��� =��(�)�Y�2��3�@�-�	�����-�aG�B�W�9I�k�j�ȋ�f|�aP�yȈ�=5�^�{��F��Ê�4C5�eN��6�I�5�d�OEȝ���U���'0_vbA�� �}3��o����������S�;����0T�OMz�F4% (gE�(QH�Sg�Tx�
�髄G7�j���$
I��7�]M9<����0���N�8p�qcOmV�Af�����b�_�̯�ɇ�(b<������������h��=�JsL��oާ
�͖ӣPyo�G	_^�]���,�� G�)�~*R��Մ"6�3lt�"�9�6wuQ�b ��,m򪺪�K���G�8D�B��"7�S]��K@��	��
���}ɇ�x�:|o�����:
��$6�օ�H)���e����.�
]9_�FaGUu&�#���Y���9�'�<��A=��6K5[�#�1An��埶��5(��wc�tV��D����f��HB��Z��.<��dZӋ?2ڑ�#tL�ӗ�L�����_i)��{�vq�Z����7����.q���m����S~���m�g�_�G��
�4���'N�\核�).���R5�pQ	8�:�!�����12 �@��T�)���^:��E����v�K�>S>o�xn��9!�7�j��L�����|��Hdx��+ho���ʀ��(�1�ȵB��I�(�b�Vkx�o�.y �X�;Ya� ����>��3�'=PeWN�c+��KqIn��f=A7
eEƯ$g������$ϙ����0 �ºF�ұ�i�J㎟�Es��P�e��g��B�N��z��~���.-��B{}&y�K���]Ē�)�Y���S9�x�թ�7k[���U��-j��sKE��`��LI��_�g�(���͂�-ƊK����V!�a��QJ<0��e���aN���(����Ld��]�C0͌�bh����TJ������e�C�o����O���"�����j�M��u����b"aﮞ�EP�@���&1�e ����a�>@bF��K�3���?H�̏s��~ 2����^vUb��c� ���uX5��㪐]��B����>�`#��a����v
�
���4�N^��RXK�)?���g'�����5��szZ/���9Y �V���/���kYj�d���z���������T�<i�M�n�9ԝ��s���� ����Dh�U��y������U4?�������t,���G�;Ʈ�3����R���i�Q�7S
"�67A�O��G훫�
2�X���r�6����ث������K��9լr�n�O,�A�мfԌ5{�Q��?f/�a�L���k�?�����^�� �D�$�0ځ	^|ӕ�Y�/a���5:=f&��^D�J:��K0x��A���"�T�
��8M�p��F!D�Ϟ��Ko�%��s�H�����uOO8��X2�$LP� �^�F� c:��ǄG&i�%�����0\�1я=�D7�x�_c4	���CW����F[r�]N�����hdZ���1�����jvE�Zȿ]<��w8���:���U�B��R��)3� ��)y�{�ad�q>�d{`*�{5�����ut8��qoݦ_�(9W�{�̒�W���39<� ª�c� 8eƦB�sb�0�|���-���C�ExK�����~_gkۭ�ʉ�|,�*��_g�Ӱ�_j�xSx��J����'v�nY�C��8i��Ak,�^����ACq��.PL���>�#��������G�T&n���~g{ǯ��Ѩn�Ğ6�����#��	f}ۘnk�a�(\���S:�y4���;6�����x�A�7d��x��GKZ���
�E���b.�8EfEt���"S��$�ZB�{&��P�s] ��z�za\b�z�E���y����M9"ZP�_<� ͖r��(�-M������� P�J��C������;PC�%�N-lՍR���-��O3�(g�!������橂�K;��E��|�j=��g�C��	r��R�����-ݫ��U6·@`6�?�g���E��	�_��r����t����߿�Ǩ+��-��uS����1��O_Jg
�g�G[T~�}�β�O\���2��Q��N�UT�%��lf%���*0�N�P�Neg���E�p)�������}�b6[��ɢ[��8���V=w���SxdE�������i��z���_#�#���E;���ao���y������%�7��|�3Ǚ��+�&��54�]��X��ٽẚ�7ٶ�ݗ�ѹ�A�����ڪKb".�dޤȎ�X[�W�u�AK�R)G�F1�i�|	�<}u ��r�$�{o�ǒ��Q?]V*qX,�������I������e��ƣй׫�-Y���?�.�����������Uíe��z�m�bݤ��a42%�j�"�h���o��4C�}��:m��1��q�l���6�|C�����rt*�C�,�2PSl�����f>/��@uT�K����?���t�d9�(��'���>R��0#����/l�S�2��l�HFHsy���y?� ��2)��x)�єUi�cP���,��ҀȎ q�EU� O�D��h��Q���ꕉ3�2KX<�8���q��O � ����K^�JV�e������Rͩ�g	��DE;y���`M���$�E�K;�� rި�M_�.UO�1��L8�~El���7�{��OR�i��� C�9m 4�����K�	�]KA�Gb�8�#��0�y��v��T@��J�#��� �<��i��A��Hʓ���?�y�ȞIӤ���|靄�놷:�DlP��/[8��I6z!��;p0%�x( �7.�� ŭ+����B���E�y}�n8�D��I�f��_���3�eřK8����H��K��{ީ���EצBX{�9xU֊����X�E{�c�Ő��� �dd��38 4�O�4�jD|'E|xYw��ZՈ�9�X9Ue�IL��,��Y��&oyj��ܽ��ɻ�gu=������5�__�,I�]��P?j����.�n0�byf����|R��Y�]�;J���]JR��2�WnWY���7s lɬD!1̥��+��]ݱ^����|j��	�q�w�3�X�ǟJ`k٩*3!!���=ި�?}���"'��; �B�u��&Ҥ
�fgO�L�	��r�M�� %o�Q�,�[��c߉B�#�Y���cn�:Ck�}��˵̀�o!ūz��r�������&��k|�4=(��̭]Ge�dl-��N���/�(&��ש�I-�Rs��P��L�C7�6�ݾ�p�M	kb�'�y����9����~�I�~S��4����l$��'�h3om�t�"��A>�3��Ŷ��*�%[������xڝ-���ǟ���mяHsŨ��0�m�\��|Y��[bajN-pl.��5��u�|Cp���~�uX�WocZG�)�/U���P�$)9`4�"�`�c ^�����o|��/��s��ᙃt�ׄR���9���^ޕ	���@˒Aq��p!�ʋ�7=sHH1��"�$���(<������	��-߁�,�����5t_�[r�&��ݦj�uD�J��+�Z�g�(�F���pT��I��'A9�&.�ǃ�]H�N�s%
B��\�Z�b@���c>Ȥ�A�a눃�ʌ�Ra��2&Y 9�^�TXk�+��f+���p8�{֎�Uk:3H�k�zć�
M��6���������{,��@k���%�+sC�����U�������b������WfI���.��!�w��S�P|w�?���9��?VUkI�(�T.��H���8"c8K���ѭ�o�r��čب�Nb EV���ܻ��^r��	ʮ%~4�<`��#�dF�[�s�L�ew���ݪ�"[J��5h�Թ��I��)*�����?H}B��h5� �j�ⵣu�yQs'fB�+��@Wkx��Z�)��ֺ ��s�'
r���1��)��m���5Ȓ�जͤ��� �a- ����?8$����X�~2f��j��4��S^��q��ؼڧ�ܤ�%����t�j����]�HO��d2��Y��-P���� .]]��	����l_(���	j�)�۹�p0:����]�M�����&�J�[�i٥��
)�N�H��PO�Hec��R�����BA�8���s�B5�`�|G�Rq�����9�#�%����ۃ���={tu�fo�]����Y{b�~O����b� l��M5��O��Ϝ��B�<t�S��i'�.��=�����r\�R&w��]<�wj��� !�G(����Q_��U �.�^"f/p�Jbeb���'@g�@B��(�1z�7�"q��, \��ݽ:O����5��˦wX�>Rڋ��#T�o���CY�m)b}m��6_y%D������;���[�ߊ����Ajk�X'�!�������5AT�F�1�"K��fb\��NW�`��.��)JNm�"~.:�`�����#iw�X�L�TC��u��aϢ��H�ʁ��Ժ�l���y�V>�)�H��Z�V��\a���k@=���84��w��`Ncێ�)�S�d��_El�H�'�~���J]��Z���Z��uĂ�g�wW���A�NVI��&�N��	�B�#�tӜ���Q �cvS99 �B�����|&8�5��X�r����aa�Z�զ��Cb�n\&:u�@X~�$��E����͑���A���V�ߟ au�� ��i�ܩ���xp�;I��n���J��Ū��adF�#�'i3lw񺉪�1�x7W�b�tP��nB��	��+)��X�����@T����2��{�4��/6rS��c��E�p?�E(H �j�Ż[R�����D�Z��
��������r��g�3F����}�%�]Atk)n�٠��0�8�%�3}�s�
�����Wq��|PPCw2K ����j���?1n<�}(Y�>�k;ݚ��_��w�����BՏ��= �� �inb';�/�Z���~�k(+��*
N6���}3��q���|�������� ��s�d�GҘc4a����a\h3y���8B6�'bƯ$�F��#C��7vvwJ����t"�ɼ{:薜��y=*����	?わ��q��ў�O`��!�L��ɛ��`M`�^�`L撒H�<�G�b�<c�J7�h��<z�B��E�P��)�<����TEc`��Y_@Á	�.�!�t�?H�
~U�^�ȉ�����,8�(���z���)9pA�M�t�y��/�tWi�w_?�꽝4�h7D��j�ܼ��U��L�sp0���J���ەi�MX�z��=��x�u�0�/���j��`꠯Q��"����l�����U7"�Vq����03>K�0C.��cz:�T��J��w|8{��4K\ˢ����/�xls�-�ѝY�Y�e�>���;�̝��>*�sY�x��?���:�E�)��I��Im &�@�3��te�Olt(�h�V]/�$�����~1�^�wb&@��]0X7��/oGsN��#p`�s��`��!�V�w��b�D�'��1��NV3y4����{�Gb
#��o0��:�������1:Y��E���vih��s~�9Q�G�sӇG\��p�QY\q�HZ����C3�s��[q��â\4�����=�&�~"��z���^�S~XGU%�4	�jvF'�M��B��$�~_E����5�B�y|Q�Le�6�3Y����H���;����-��ϟn��?�9�75P뛰���ޣzp����(���7���uT�'oo��J��ܒ���^�J|�u���a80��J0N�f���n��(Td�$�-����������I���i�0����\@ە�̝Y�l��H�y3�ANX���y�=B<��[3d�f\���B@5����e��FL�e��V�Z`��7R�Fpl���ϒ��f���4ѷ7h*���~�RO��Ds���>�.�$����á���%[,Y���Zb�u��X��h�z4����H���{�pU�t��W��]!�� �`����;��x����($Oj �f�����'�h'�3|sh��_v����7G��p?�ob���V�d�T�o�͒	�-~ҥ��w��#[Ç����#n����#�H�n��s���I�1V����I��*R@5ͮ�V�"�)`M�Z����D�� =��-.�x��ȫp�h��D�Z�U��%�����s"���N��H=�s�4�3s᡻��ۓFt,<n�� >�r�5 > &wИ�3Mh��=���|��'�k#��&S���G��DN�n�����5%�g�F�[\�J;Hg�z�8S��8p���Ν�*'R�{�F�(+�A����|���2Q]Z�|���������\�g��7�i+,1g�Q�\gokǖ"�H_�-M�20��4�h��I�D*�v.!nt�j�,\����qMi�ҩ�a���	�� 
�s��Iu�.��i$��6���M�ԅ�$M�
�GR>��QM/տ�6�Щ�� ��`i����f�/R���o~тE+�߈���cOxy/] ȝ��4���(1zd\W���$�K��/\��It��1�W��pN�2{��cn@��҃+�U�-�E,	�ݹ��
qӏ*(�~1���dc���e߶:v'�w�"��J�����c��K�ǲ�DHQ�9LFvu�>'j����G�d@Jo�t�+���F1���:48��णb0A0�gy���5%����g�z֢~���^9�A��u����>��]^�w� Tw�W30a��㯜̼䪁p?"yB�c��'(�qޭ	��z( Ԕ���}΋b�d�m�4OL,Q���E����jY�X�~P���e�d9�pD��7�"��D���JsFf��^�;��xq�܊0�=	����0H6G��rz�$�7���6��WͼV3;	�Un~�Nq�Ol*=~���Zۯ�_�	����Q�H��.58�
�o0xI����Z�u��|>��������||��9�~7��=�F��<d´�U�BR�X�oMXn��l,9�l��9��7ea�����@��(+�"g�Tgt�Α�C��v)�#���Z�3;� ?�'���ƳMoA�DZ�h��>��w1$�����"��SF�������@+��L����;�[��YQli}싎�;-����>i���3�	'��I �*w��ZA�=:���Z��/���3ĳ7�1�mq���T7c+��K�����b/c�ҭ�0$����WH("e�.e�������~�:����Aƿ�R+�a�7�}fa���@)y������G/�u�3kC �T{K$��B����V�D'���)�����u?�Q'!2�^!XF@����n!+�a#�T�MF���4-��G��`��2��~�-7�K��j�Ц�r�vc�P���>΂x��U���.���[�<�,Pήt1��//����x�'�A:��m�����ϊ���JH[}~��\!��EoD����s�J_��͈��T��-�)hQJ:ʱ�ƈ�MM�T�p���$�T��3�r��*�����ʨm�9
n.T�WT�QA`�Y]	�<Dׯl�\E�)�
�T2��-��^�I_7}O�*�~D�7�gH��1��Y�7��ǆa���O�n1��Ⱦ���3V��1$q���/�i�[K���%�f���ZF[w��X�C�Z�޹�9���ǵ]o<�F�>�i��mv��r��>5� ��������S��fL����Od�	r.����O�BG�?<#9X��ɮ�Eo/l�o-D���&�B�7��h;�)����@E�A;[���(5wbH_�'Q����}؈�ډ�x1<p uH���f2�R��˥��f)#Ђ�����ÔRteYn�$\�T���wX:)@쒏��Cj��sL�	-�_��i��I	Gԭ����Ѻf�y \b��Bq��S4��~�~���gJ�Gj�Qt���?�������������_�*��v�JܼH�P��� �U;U�e��,R��͎��0]�����0�Z�҉Ж�9��6K��a�׎�c��s��:��\=��vr�����gY�%ż5������0HxX�1�bߣ�5̸EL�)j o5�\�Lb�1�(�o}Y��;<���@ߦ���l��3z��O�HabC%��I�S-P�f��?:��I���;�R�Rj� ��H\�j�/��5�ɂ|�U��W�O�� ��i��)�H�d�{�w�������yx�Z���i����۾3��N�>�dqI��xs����I��N�	X�r���@'F"�
�h�J��؅ƽ���\#�MEQ�bl�;x��oA��i��̲�V���y�.�'�1gC1?��ȏl�G#;���9aOb��߇;#�����s�C�7�v� }��¸U��E"���@	zJpwg��9�)�ޥ\~�kf�л�2'ƞ�=]Q�>�e3_hI�>TܢZ�ި	���E#�bb�l�\�.��@�he��K]��pa����M��]��ů��6nռ���h+-�&�Չ�n�����T�uu�[]�`P4w�	��(�윹�(��$����T�d�N��e�:ì��f⣚PӃ�SX[��11�x�}J�pߵ����Z��J��s:�QE�T�	оK_�����q���6
���n��e��F*�@����ѹ�Go��"�fwu!�"�f��SjRH��?���ob�}���#�
�qps�
�2��s��e��eއ��6�m"C8�v�;f�?�&k�����#� &��h a�qR�.��
�b���M���ک��Bn�#:��N̱�_���<RT��(UC�d��S8���w?E���w�^^�xA���J�к_�����[��gW)_߀4����
ԋpA"0��m
z�[ �.�X,��6�E ?Qd^:�C>C�V���恹��3�������k�_�i+M\���Y������L���A�v|xܿ-��Q%�\��>q��(2�?'�T��,L~�C�hc��1"���2j�j�ɘ��l���7�u{�,��	� �[��l���E�{:.Hz�����M���J�y�.��Z4�����x\���g=a�e��1$M۵�Z
=�1�=(I�Ӫ��F�õ��
�ppn���H��f_�Z��u�Hn�r�ɂa�h�B��@{���2���U���<����Z���~`(��AN�@�M�Z>�,�D�}���
�DԘb$s�I��P�-�]�G|3���Q�' �)RJ]���s�+g��$�J�!I k2�"��\\#%N�D�̤��P��U�Ǝ7�ߨ����Lh��l\�h޴�!� �o���n@�
�D� iVǕ���p%ѱ��1�`��� O
5o��!2�������e��C|���,����%�킯����z��U��A8ʽ�h�c���r�(�f�S�]e���h�> "N�l�&�}QCw�Zz�齛5o��ط;��� ?�>�q��TFx�g��s(�o ј%��C�5�۝�BxKa�����P_%�6�f����d�y���|��Y�:��[��Ex�+~�Oj��L��S�`_��y�J*7��hɲwC�x�_��*��8��Đe8%��4�����t`���	?������I-ّ|��.��,yȝő:�V�� ̵�i���Q���r���E�T�n�9K���^Q��L ��j`�r���]]���5�%&5��EWf���/z��W�����'��.��%ꍈ�A+\��]r^�Y+��fk���� 2=�`\��_���0΂��� {��ZU����~�����J�?�*�Q�MOB�3�YX,�`q,H�:���|X��f�lv�eT���oE����/ˢU�c���&5�T�xP�հ���,s��5N5��Kw���۔�練���V���ބ&ϣc�����P���̞$#M��.�|�,��^�@%���6�k]cL�^i���%!5Vx�������i�|\ ��}�H͕�ǠЧT�~_���D�*uy\��6pV���bGܗ߇$�z��qt�}|��J��c�W����ZV3!��=f _Ż��3l�C��J?`�ֺ�w| ���"v�>5��X���-v5|7��1Č��}��'Ə\�-���H�<�@�X��񌎦5�'U��Z�D�r�;hk��/ڡLD�Ů�k
�x��Ga���V�3fg?�:�����u��V��������w�h����_,&p�Αu���@��f��X�S#�FV����`����~�z*j&�i �LH�$�3�
n#Fu�ƾ��d��<�,��1���o�����	�VV�W>��{�����f�hv���!���?=�v���|�j�M'�
��X��'��g(��u���ڜ���B�8��=��-�+��jv][f���N_[�m�~ܦ��X�Ig�1�kp��S
�d����˟�Ag�y�t���B���V��@�dAj&6��7�m����q������_/��﷪��t>��<����u�i�m��/V-�[1H�ӚD�����"$�L�S���j\�kj�Y��x��َ<k������E[C�C�x@���t;@�+�[��I�0Tì�G��m�Yۊ��>34�2�e?�/�B���N��A(z�>�I�5Aܜ��Ҽ���Ş���*�����(3�B9�΀�|K'�ESʰY�Z�����N�@�v	��H�Pm.�e�P��E	]H���EK��^�:\��ي����{˄��Oy�;y����u}�A���Lȿ�Dw0`�4�B*2(��!�@3ؑ�-��L��A�`H"�qc?$=�Ć�+/��y�x�~�O�L�ԅ�/�1\ֆ˒RcsƝc���5�#��4��)�����|09�m��.C
se	�̳I��&$�z��I8q�Y2�䱼C����^r�EWL��=㷨]���hd�QNc�_���\@����������\�K�U�E���L�w��d��o���гJ������`)N�̶���9�E��yC	�-B
���Ӡ8�`��GV�r<`��-�q0[���Ҹ�u� �R�w�Q�Ȟ��� ���5
M��_�­����p:��y�u�}�92�>��g�z}&ːp$��]ʦ����G��9�g��u�$�r݅��0���[�۠5Rs��Nzў�E�)R-��m�bqp�r�ʨ~���U肀Y������D���Î�o"�YINw�uMF@���'�X�ր��߿��Ex/���fX�6����ż\�TZҾM�X���(@�vP+\�W'Yg�����L�*ق�.=Gcױ)w�L��C~���k��y�i�X�Afn+ћ|�g����X�	�_����'�߲i@�o��m����uTjNKa��/:�[2 �q��Q6L�ZDilrS�u�S����oy(�P�NIGg�؄��㲭sIwe�j@?Z��z�.B���I�Ѐ�+��z�|϶p�E��1fL�Ew�W�l5�{������=�$����E��%��f	�Mi�صG*v������o$��z8�?0�\�f���E����v\T3�WW�$̬V��r���?�&�����E_wo|G����=X��@B���Ϭ&�b�!R<&�N5ħ�]%V�`ky-�+U(ZƂT?Z�|���3�wކ��Eد�=��F�!dX��y�<ח�=��nX~xQJ�	4ИI`��$�.���J�^�Q�[�G�Ԯ�~�3������Go�;1N��	F� Z�=��Z:�[�~�>>�eȿ�?���eһ�4no4[����̊�,��R2�����,^DF�b�6�*$�1�y|S=Ȑ�
Cm��1͇e,V{�[��T��#Q:m�a�:E�n	��BQ����kxr��:���a ������H��M�0���媺���!ԯD:i�]�myiՄአބ$�@������h��Q�u�p}jO%�TX����0��̇�����0�������=�u<�?IM�Dd��H�X�l*��?�N'��I�V����jq8�xS\2��p��g��xfl^�PŊ��U��)gK�j~8�֕�	�ŗHb�'!���C;[�B-��kz��C��6Xҿ� 'ܚ�OV���B��y�l7Y��8�B�]�Xo*{�`�?��?�����܈<�/��`?==�������F&#�i�]c^&���%��Y�Qh �q"�+-\f�Nkdɜ�ݧ�>�����NS Ei:��O7����L��&�O25v�����3���A̻OjQ�R t�����B����5$�Jq����������~����	Sba��f�S�9~q�J�V-�z���l����z��� BW�s�5��A}�.�Χ �3��)�
��`��gs/�>�Co��hj���R��Ȫ�#8�aWn1�=�lD��Ӻh���>L
��?�~[�Wd)����.`v��!D�$���Ъ3B��@Y���r8�^7����_�@��̬�R��L�0�F����Vƥ>�K��y�&tJ��`ʙC� '�g��ma[}+9@֗'Ya�1ٜM��ȡO^�A������P4G̦��0�*�@W�����\ti�`��ܱ�X)�[��u�jɋu$0�q]#�ad<�9�b��6��)<=Q�Vǈ��!�Q<y&S�|�%�u�,�����&����<o!\���
���J��<F)��EMlH,�`+�2n�Ċ�����z'��>n��z�܌���3E��P�-�*lV�f�8�������}ʹ���d�^�Ӏ
�ԓ���Ŷ��2�
e�|',�ѱcM��z��&q�yY��i���*���j����
��dL���10��C��]�j�f�	��dW�Tqwf�����;��_��IJb�����l��f���[k��_�V5�X#i��j�#���m	/�$Ì�.0	e`Z�NtQ��μ�����1Y���UG'�a�*nxԃ%�Hm������	ݟ�Ȋ�ב�s�nėh#��"1�Iv��nw������X+�j�t���t-v
�����fp�����ĳ��
��_�
�y3+�w[N�A�x������$)�q�zfua>�>��~ֆB�;	Q��!�ɫ�`:�
��%�FX)��ӈO& [�����=��Y\r��v*�H�h	����,�l����ם7f ��+��*ޗ����L���-� ���F_PRB�i`-gyad���u+���orK]R�������
j���y�oFK[�D��z*���&x33ȄJ8���= 6��[:^B�5b��7�,���2�;?ElP�����/��ќ�6�ש<�x�`��j�,����=H�s?єu-l��x�y6_�+J�Qۤ��<�ʔ�Β���U��B��x��������ºo�4����0�`$��p�=s[_O:W!��|����<� nn{=k��y٭N�B_UW�x
�Z�y��[�P�:�x`����Wrꟶ�e��ys��0����]}��O$ev�����!�R!	�����@'m���lW��'���}t�3:��U��$�,�D��q=8�s�r��)������L��-�?����9h������5��8�c��/�/s��]���wo$�2�X�ҥ� �MD��QĺeC���d�0�J����j#-��N�����9�x�FӦ��L�82�U)��)�~��w�c����ƈ���G�]�9j^�FbG3��H �����R��M6��#�5��SӪ�  �Hhn��xO-��xT�b[/�ܟ K�������N��l�O (��tBJt�
��e}ԧ�����(�I!��&)�e��dJ��}K�J���vL`���1}7�<�GKt��E�)�t���e�؊?ZH!�Z����4����w�����A�b*5X�x��?���)|[�
�+������l��7d�_)Z��c���g,�Ҍ����I�{�����4��uD,^�.��-:��\��*B�����X�侓�y�YK)��)/HF�yN���8�$��#�i:�%`���W�e6�r�o�ɷ�8�/��s�^�:8R�u�c��q�'>�r�vÃ?��r�3�6}F�Ru�@aI�#KV���E���t#yp�
��c�@��<����������'\�xj�ul�㑗=�L60��~m�iN��.O�C��h��Ήvyʸ�O��#n��{��mi�~�~�[9včq���kLp��j�*�;�&7� �F���������&eM���D��Y�ӿ~o��M�q/$���7�ڣ��22�]�8�
��0��+�n�Q�f��J��sC���j�h�8sZ� �5⵭u|%L{|~nc
A\��/ϴ�M[�ͺ@M-xk�R1����x���`��}���&t�2|��n�Ѱ3
�}O�S5b֦B�arq՜RD�����	�~�OT��ӂN$m��U �ݖ
�L���{ȊE�X���1��T�1:�=qR�Ժ�`�vk'�޾�a��Xt����H�=w֦W=ڲ�%PǤ��u�6�ʤ����5�\v쩞��al�ea(�s!K%1�����ymf�+U0�)W���(�aH'A'�2,MV���F���,�rn��U�6�[;_�9��i�������mld�OGԭ�nTt{t ���% ��q ���$�L?J�`ү��%��U�k뛻Di%v�����{����qu��w��7�ꗟ�ˠ�N��?�}����PDM����3;�]�Klj�o�Ia����0qSF
�ԕ�����\�9 ��y=���������٬dn�����H����fc�>0(I� ����K����C� �Z�Q ��r���:���^�('�)�9��c��6�l���"�$���gE�j8sh+���U�]g=XA��2�`�����D���nL�E�{��!1��~���&k�@0n��H����aT��$�����GS�� ����V��fq��_�_`OA���ħ���gٌ�vc��SPZ��!���|�C�!jʦ@�CTY�&�܈�`��� .v�R{� �>>u�i�f:�nϺ�F3��5�c}K���l?�g[#�_m]�$2:�[�tK �,Kx+���w����{i�ͭ�GI�%� ��w�_�-h2�&M�&Z��ԗ��E�A9uI�H�)l[��	��VjY��5��~�����{DQ��@ߢ�������>r�	���H��吣	Q\�{[3��ǡ�%�L�_G�	}�Jv�qd1�f�e�$�0w?�X�r0}��=l����uF�K4�� �)����m��;�*�"=��0�ܙ� �Eb�r�l銩�h�T���A�3��/̣�g��\�뤉)������NEsHr��A�:��?�@�5����]KT�t�@t��l!�Vnp�2X����_ᨺ,v��kdt֡��X4���3þ����R8�_E�±���]1U�%M�1��������m|`�'���{��E��f.���9��k���q����J�#�3M��N�o(<�G����hk�_%c2�R�X��4��q�
�=�瞠��J�Y-�Ə�X��ڼhN���6�@'�Zޣb���:$��\m��6�A9�cj���kK��[Z�b���Y�ƒ7f%����$
[�v$��wB��!�vq�:ئ��/��k�����|�a
�%���Ը8�]7�X)�h��c7|�Οoҭ��b����f�8ীȝD�����M����/�%�n@>��H��"�q�Y\�ra�2���غw씏1���l��&�'.KvPA��nm[p<J��h4X������O���l��a�6A<;p��߀)RE�&<1n(�㜡�9<J�1�/V{L���L=~qa#Ю�Uy�Yq���,���J����
���?=�~J��"�y�%�"���g���jd�֠�3[���j(���P�B¹�ia@n\!�l�R�6kP����K�IAz��?�2�z^�ȷ"��,���+S�N�\���2x�<+ќ9װn�h�_�/�E3����d����"�]�Lm�^�wO�E�3�x���[�?s-8�PĒ���l�bː�J��EdgS����q�,�eξ�2kUF�©�,���f�K6�h��ͅ��z�e*���Zd����i��*�}���7���?}�n(�`i��N�KtN�����NQ���
`}(�<��I��Y�����<�Q��:
���&��#��v((\^���� 4���!���w(�ĩd˙�������;R�{_�j�������C�T���m�����@���En:@5l�k{ta#<Mu�ig�r�����ʱ2�XHtꪝ0͚�d=���LIt����H�<d
�nh�ms�jPn�r� ��B��L�9����<�$��b\�e��i(��pn;K���R�ԟiI���mEE洙����(���t��	U3�Hlx�<�	//�C��5�/�A��C>�fl�b�I�ْAM ����8�
��so�6�$�m��
��i����'���[�L�\)&\
��pd�ON������Y��Qq���/C�u�#`jU�z���ɉY�3|��c��i3�v���Y���f7��&��h�M�:��|�Y���'��j^ߤ:3�?����:-�(x��'��5�fY���Sߕs
��z~�#}�1���<�4�ߜ�oY�E���#3Z���D7���|���Y���S�����eKB�X���lr~�����oqv�H9�z���ɤ�~b��MR5�W����j���F�д�����.���qtֺ�S�*�ZaӔo�l��jp�: (jJIyz�I�0r�9W�<X��h#$� }�31�iҮ�K;�0�B�S�=ϗ�/�sW�+�wHjb��K���`y6�D�YڌY�P�:E�*�T��W{�<��N��厃�e�Q�w��/3����W�rFM��'�H�s���68�A�GFy@~y�2����KN�_.�PX@/ͤltꌪdߦa�n�P?�P�ֆ,�D#ښӍ^���o�,��<}�w@�y��{���˟�����y����l�/dŧ��YE��b��ΐV�gwEns�������l��a������~>�ve��E��x�Ĕ�t�*�NFI�bNHh(�G��Z|�0��Y_XL8���yG/�o;�C��;�#��A�p�V$�%��	.�j=;�5�԰�1��3d��.AʷY�@�\l5�y_U���M�?	�	�#�;��� S0J�z�P�������|%V>�,���5o�]䑖p3��p��+6�(=�DM��ma�q"򕻛J'������4�L��� ����ca�xZ�@�_���u�@�2�ص)��o5F�OF23���T�'cq���C=;f�zC��"s�����yjq&��zf�ا�@��1C�;�,��f
BІ
p����$8�vk[����1<0(>>���+m�O-�~�_!�ń�^�Hٺ�t�.��� ���lh�u��1�����-(h�4�b��F���N�?�yR�
��X�>�
�?��vHv��̞��lN=�Gl��*��dyK 	��K�ef0���p"�$�+B5��Y3�cJ�,�~�*n�NQP��卟+Ji���l�KN�����gg-��=	W��94�"(̨	<8���\�z�&.!0��H��z�f�"�8w\��Ͷ`�[���=b2.�����+`�wi���Q��f=�@H"���f������_��S~���4��twy��<�� �;��e'O	��3�e
�Ό�ۼYbI#�^�B*���'��x�;�F�֑�m,�"�_2��z�7�94Cx�/�?d��S�Z�zz��}�U�n����k�W�b����� K�= ���H7�\P�(��$NG����)&�������!.��]0��=�Wt�I��|�M*p����������f�wRL.C�K�WU�X�r� �,�LTp�G�LO���.�m��
(��|UZ)p�z����s�d�C�s�=��<�eR����vh��R���D�H}�k`��1�ŭ���<��Ҥ[0O{\(�b�L U�~L�e)�A��e��<����B&�Ԛr��m4;w9�����j94"[Y�@����	��������6�hY$5�������e'F�����Mуx7N�]y\�%Z(-g��折2���!ȃJ��z[�ఖ�JR�Ji�G'�����$��~C�M+b�i�IV@O��\��N-��� sNFgҿBEʹ��봳�OM�Ѵk\Hظ:_<�g�s"��Y�Z���ӈe|���;+]$s2���\���!�V||�� o���n�ӾiK��E��&�/s+"<�|^��-z\pG���MhX�&�}[Óq._�9(�����E�o������(��y$��]G���[�����`{`����/�\��	c�����Ԯ$�]1��i���TϹ�f>�
嫋����x��[|�����(L�� =����!�I׏����me�^�ヱ�j�L��tQ��P�)����$1�R��)�:+ݽO��U*���>=5�n�M� ���������Q��֨���1⾗�!�A�"H��":�C��;.e��r�ʶ2�)���4C����z�����CQ�M�IU��(1����_ 18!��rT~�ߜ	�b�ǵ�����8�<�[/|j%��~|z��wJrqn�J���������2zժT.y?����E�����29����V�9�Cm�W�z ţ�~��%���Ť>�5�7[\[���oe�0˧=(m:��'�/���6��
���2�h�ݲ�%"���f�pB�H��4�í5̗�,��0# ʹ�$�*���HBP��P�N'����'��?�]�q����@Lͦ�W�fǯ)��Q�\�ظ������m��f&j�݈B{�}=��D%j�V�Aנ����:u��=5��V����Ϭrߤf�C��5��~NԚXV�|�,��x�"
���l�/2hjK94[gQ�o;(!|�ŝ���Ws65�7zۦ{hB�}$���˨!�)�L�$���H���%Ű�@fǏ��өU������*��^�ʺ���_�"��$��ϡ])�jE����A�C�폀�JK#)r���h��@W�-&ǲN��������mw���� �Z�^���"9�!5�S���0��\^U{�����a�C?�M�p���ə����nB]��½s��|st�ù���5p&�' [:�Je�s���_��6o��}�r~@�<��{�(tV#5\���!Ȝ�@���B��C���mR��T�((Qmf��Nz�	�����b��|<e�������v�s��K ��� GH���=h�����0�h���"#\�8�Q^8��g�S�M�먎���0I�h0���r9>�;��i(�=��`��c4�ǲ%pӄ�����+)uQ8n:3|8+T���5Χ�Y���2�V��6J蜹+ՂdJ�� q�W��/��E��3�Y}����C4�C���#��U �|H�|:)>`�;��f~&-GI�:aR���$�&��=�!�,�&�H?_Q0��/�V6��/��.��	�U�>�}�&Y��&dN��FN�mB�~�b�6��ڑQ;��IE�1�����ئ�Mx9��.C��p�Џ��7	�X�B>eR��0V��>�8���
�=��_
��Q�p���{'��_r������(�v�l�L  �G�c^zu�V컜$�A ��܎~�w��|��^���<eK�s���ԯQ�/���y�"���r�9/�[ �t��� aD�f�"��E��!�ً����6�>�����ɴ��Aᕆ�z�V�E�s5L��Y����L�h�PZ��Z�k/��bZ���<��8W�e��-�pB	�	��4C��(��r4b�h�P=�B�C�=x�!>���6�˛s6Ff������ޟ�����v��4vh���$V�0`r�@c��l\�q	&�'U�|�k[>����)D\V~;��\�dŁ'��y���i8F��CcH�k$e��"�O�]%,,�L�D�z��4~=��rX}��>�~m�͘��M�z����Vͤ�FRA�&bԾ�T׻����V�)�:�-�z���k1�#EY��H*�z�33�YQxh
Lq)��!9���yѱ`ɓu��W5�8{3.c��eF�F/����[>�NH�% �9z��X ���N�e���C����~��{j������eaQ�iXy���	n��Q�?�+˧Z�Y%�F�#{໯�kOZf����c��CΗ8X.��g�8T-�����5�i'7UYX3V\^Ķ��^���$n�A>.�EutR��2F�6D��}1�i���B���^�e��M�.��)�.��3�%�v���-k7������?h��0� ��?� �DC8�":h�S�R�&���mfq�j���c�?
��@!cI��NY��=�; ��4�Y91޹��"{���q�_Z����e E��X�	��K�C��>>�.�a�* ��>�M8����8T=��=aݠ��K�`�PHP�ڰ�h�-ǪU�1��t�\�(�.���<��p�7�F�<c)���L��!$`��R�6��� ��o$A:H��l����zQ���_�CI�c�/Ϡ�}*�?���/��O���u�F&0ø5y����4lw��W�t�W�	.�&h�������g������6&v4B���r
�8��5N�ѱ�W5���\�#�AК
I'C������St��ϳkC~��I��1=�_fE����k]��=��\jEZ�#5�T�ސ�ėZZ�l����)��n�&эnF�		t/ʖT���lyR�Y�\+U׬�-��e&ŵ3���W��{���~�N ��{������Wۧ��#��@EJgA-ܑ�eᅦ3��\	����n���L��.��I�a۫fkv&	� ���|��ש-\ۉ[��PLͥ�$x���b6��ld���2'��&�������Rģb���l��s}����z%��2n�Z�ۀ�C	�T�����|�Qfݗ��*�)ڐ|):�]�����N������Te�����j�l�d*�s���m��J�q꾋Tx%w�wC�m.qZfH���y�{��Ds������LcQ�z	T������'ã� ���ܠm\�0>.�6IP�W�xS��+�8�-W����,��+9�����%�h<�=o���C�v�'Zw<Q���m/M[.ޝ�5���h�LbL�� (���[Ά�㠆�g6ny>�Z����&�%֔4��i�~��Y���{6 ��P���tt<��T~�����Ev{�a8�21�>�����H��=�o[]�a��3�Lg
�m^��(�byoN#����{�+�=�u
9�́�ǕW�.�¤�0�.�M���^����GFx��	ުe].��R�����Ĩq���u���9�ytC�$�"�)=�4��ِ7|�W�r[�\��:�u�d�b��|s����{����sݔaڅ4uH8�՚���:��'�0�������z}�^�IkuiB�l�U��I����IYs�|2�z���wTGxA�L�&�E�������+�����\{8����GjÆ��nQ�Qy#��ID�t�����0�80�#�αܥ���N�� ^azF��'��O�L���=7X�Toi-��%eG�SF�Ӿ@i�R��L���������i󖮚kOD��Yh��S��O�ocC'���>%G�>3^˹��H�q��Ss-��I���1�Y�����sFY�s�Z�y�w�{���jC]4�U]��?1�`gl�:e<�5��4
R�<R�5:�T����}��Xnm�P�A����SZDԞ�3.��(�?���N��%��~��� 9T�!n�x>�cbd��sl�օ(g�%=ى9�c��|D��7� q��S4�c�Rk�T���5!�a�Fw+��P�# �\<=ۓn*�O�~�R��E++�l)�P:����$Z3tH��*a�V�K��p0���{���ڊ��66c�Ҙ�r�j���3"H&�0җ筑��l�t��iZ�.�)TQ��$I6#�T�3f��r��u��.�@K�	eꇇ[6��1�A�#+� ��X9�"��QB��m�8�m ,`����u����G»�v#�xy����K&�A��B����-��c�>��i�p���q��H��\���Jg�����_ra���2d
��in璲��Z��?���b�1G^L��5ؽ����Y�	�fD��*=ʹ�
+�=$	���ē>�>�j���ٽi;�����d�ߓ�{�:�|N�E�*�+�+���נ`C?N���uۦ�b�fb��$�@>���f�fw�AV�6
H��?bO�Pv������9g����3�+���|R8�)\.9��'�{?�늬���B��/���9g��>�|ҩ�c��������:Qc��g�}/8�7G~G_����\����Z�w>�G��6cu�E5;9G�����ñ���*��{�?bFJ�_-����h�!�+;��@<l�~���S�%��v�ԟ<<�\v7��0���v��R:��B}[d���`2���s���8Fw&6)&���=@:o!̃!�����8y�a����N�)��ZW%�?
�ڂ����T�H��|�QR�e����.��R�5�(>�\W9�R̓��`C;2��q�ퟡ}5j��V4K�e��7O[~�ÀEF3�UX,���^�7o��1�2T�k��{D�Ec&�_��@�Bu��K��٢�t�D[<u5ז���|��E$���]4{�F)_ks��H��9��z�,����ΰ���d.~/=S�L,8+���+���.�;���ڄ>��M�~Ft�ߌj�j��/X�L������p����Gֆ�T;���K%'�$N�&� F�,��ln��'����P��p��;T��h��2�'���W}��?Ĕe8@r)h������r҃���>���H����?Uq�\y`����c,ڀ���b����s�n20ȽOȺ�l��u�D諍�!z˘Tg)Ę��V:����Z�'��*V�X���m���D7�=f�w��s�\GP���z�\KT#�Bm�n�w�؝,qs+ƶxSR���8ȯEz�n�&~�8V�j�R���~T�o_u���AF���r% ێ�f������x�w�4���,M�G1
Ŵ+����������#>�`���T1?����U�8������h7P$��%��;$N|��g�qq�lN+���|sRCO��C˿�D�v��ӣ�*[^e�y�a7�̓���p�5��T���v���7���늈:�� ��1ll��e�wLtл�q��֥\�<2��c�����9�!��*�*G]��N��QL� N����i7s~]�/�9�vݢ��аXd�ȴ�	�IT��V��'���[ng����C/ܦd�Ou�˓eq ����x�͛:��<�������
b�o'.C����t^��	/)����_�㠒Na/�L���i�˼�P�~&��1zX$" ȫ#>���S����#�+���yB�r���hS��ʺ6 �۪:���4:�ަ��1ѝ�,�z�M��6i���6M~s1z�h�l��Ґ�D�hp(��w���18<+t���.Y�e'cc��u�ȣ�}�K�'p�2.r�7x�B�,j�:�q Y�v4�?ZˢI��(�!�xp�)�H��'+�	{�G��Mނ~$�`�R�(p�x=S�G����6�Nn�����qr�4n������|e7�B�� �-�E���q@ߧ�OomG���N��R�zW�� �����E�o�pϥ�S
ڀO<[�P�JP[A�p��1@R�}/Smy�³<�\�l��,��[cx�v	��Ϳ������z~"��
�O;A�Z�D����p���]52�e��������Qe�o���Ƭ�%���D��?���B���k-ԣ��a���ٸ��i�4�Ka7+o]Lȑ=��rfc��P�S^1GN_���_��m��Q��ʷ+���,ʞ�����8b;J�I�-��~ ��l*�R��)?���#|�y��g:,/㾍��8*� ;kx��Q�]���SLK����K�-%w�C��+lO:~�Cv"{��$�1���.&���:ET���"���鄚���[�W���u�q?{T�t[�������&U3�u���]�"֌A�vlq9���<����3#t	ծ�Yv��I�����T5�da�o���TP_Ս�t����v����=k����z��AU������~t�\��]p K S�ӖA46�T@�Sb�L��{;0>i�%�+rCR$AC���<0��O�b?��r�i��cP-�~��&��'W%�	�n#=	c��"���٧n�)�=���z,���K���g�ɴj�u�]r��!�43�N9oCR�|�XkA��}Qա�Q\}'ɱ�z��=4�_54Ċۍut,K"&]>ɒ��	���\i���!��aT��(_:�僨ȏ���F���4�=Zsb�S&x����M`�*%E���\M̀*,�B���e��]�BE�fP0�f��ح-BD�ލk@C�\t�°�h��v�'�C�����84��̳ɪK�fB�V����d�WgwJc���#_�~����ǮO�
b��H1�i^�y���x��=���j �Q�'k���F~6�V,\/Q�2�k.�d%t+ȡ)	h�+v���ߩ������Z�i�]};�5Ń�!Dt/Z�Q�&r�؆�̵�^�$3Pŉ��
-�>�?&���O6Y�A��d���K�>j�����P�T���z��8��4���������p�^�NA�3&��~����R�N�goEK2iz���Sb._h��|:���Ç��w2i4�����+�IA�lc����f��X������;�e�'N�͋Y0�T���n�Ȕ���T�H�s|���p��"��ʆ�Gy�ae�cފ�a�;�`�Wޏ*g����c�=k�C������GqBD["�D��Ӹg;��1�(�q����W;�_>��H�n�A�� S�(��q�3�-� "$����\w�� E@�CyEڐퟺ�Di�\JȄ����t��L���\����ؒyzu��ۏ���L�,��~���㓈�9̋�tߠ�m����"�L�Y�J�)���$� S'�k�$@3x2ƄY����{LZUUl���^�j��� �:�g�7K�֫E�����B����k�)�ٖY��|�S� ����y0E<�|�e����(d�c	�!�R�H����وJ̘*�6+���^0|��胍��7з��e�Fی$"{��?�}=����2��_q_w���)b�"W�������0��?'�{��RT��^�L�ɴԛS^�}�$9s��t�oύ?js�8��l�H'%����ӿ�./�L���Y���i���OϞO�����s�"*s�pa�QG]1w'��;��,�FA�˶��[#A,����2b��8�<��E�ڔ�V`X@e�8����C�gҋоp]q�'#�?	��j���Hl�����V��_Xo�u�6,�ysr{ѓ�C��;6.�Gl���Hh��}���VJ��"�ӂ�/���Zty+~�����,��%�i�L'~TtQ�Ѥ� �4��i��^�ᵫt�/hS!p�K���$�L$%���i	U�ғ6�b-���#�zUH�t��6��P��4����V}���>'Hwy�P�������:�uf��Y�u��{��
y�I�Z�3���	�o�]��2��|?��m�z����4�m��3�^n�#޽����yX�:�GI�깮pR��W�����S���q�Pv�`�np��%�����&X[4�S�?���^��Eмe@���W쏴�LJ�����"{��n+s�g���B񅯄f2��$س��\����� J�*�c*4H#p��'���|�HEtgߙ�S*��4_w����aR��P4���a4ayW�iᑧN��3y^�K�����8�\w}�w�IY��P�ȅ�BY�0ޫ6oCe@�ۊb��t����~�Y�1a&G��9+gl��Z\QCI�f������F�)�.x��`oߡ����ߑ�!�x���"��qJ~zźp'�<���r���M�v\^B�ٖ 3t��d7ٕDU�7�?3�b5W!x�q���+N;+$��o돉��D�3�`�������Ȯ���.���\�_tԣ8/a�ljh��M�{X�ݬbzx�R�ݬ�+8�r��	���M�������� �u&Z\���I�Ԉ�C5����nH�\�Ŏ6�s�i�<Qj�](_�ܺ�eg:2����kBe
J$'-�=�����cAL��ܖ��]~�^k���]5Z:�ih���!��F���nG�K�*f*Ij�r���D���u�Z�P���Pף�X��sz �v�])C\�gQ��Bnu�d���@�^��0�*�_i�D�h�-�������'�아g�c�q�&�\wF(��1G��G~�����#%d���\u3 ������$ۯ���K��3X���H�z�M��y�ŖIM�;�$\Q�f%�Gu�[8���L�~oO�����Hd����ᆗz���4 &<�����-���br���R����Ȳ��3�;4�p��f�iM�&���r�jd$�uP�^G��޸�}�.��W��nD#��)��j,��Q�V��%��J���ɂݎ1����]T�?�1�lLk�}g����W��O3"f�R�ɫ �:�=h���t��y��U3���܇���e�lR��3MX�nS�3��=��Z�5b�{����i��':Kq!�R���T,�F8���HeIY��>��-��e��y���F�8���d�}��m 5o�e�0�Ѣs��E�W-E
���v��j�7d��= =�/}�7h9����
T�(:�$ RlI�����xs�*�IS"`RXK?�>�_�� ��r�"�ܸ�|vd\�#��<\)���+�c�Џg
�	RS�S�,q��"�e,�S{�^���IM�{�6�_�.�� EǮK��ѧ��z��@	=�wX�{�ek��WM��H�d�E:�[:(�X�6��oC�?&
�.�-���Ǐ�>1P	*��h�-��=7���N\�o���
�,�EL��57��t�+�R|D�T�P����K⡶��*���dt�,����fIX���$�]M��~�d�+�U'i�8��ձ�=#�R�����8�3����iC��k�MaVf¿���db�Æu�@"pF67���2���b3A����5���v�n��%���#�J��U���|����P�����U���8��%�Q���p��붕��G�fJ�:�$��u>=Io��_�χ@�뜉�|���t�l���u'�(ʯR��q�!��M�#���9.����
8�+�mo����~5�P���QtইdZ�kD�$����1��B?����}��ʁ~׎��Z����lHA�ԶlU��#�>�i�e�K��;�f����/�/�c#.TM8|$wjݳ��P�Y(���U�m���d4�/Z�<�S��d>�Wn{���+�%�\��&��y�����vH��\�E�!��G2�^�7va]ӻ G�����Nf~|��M�����tX�<]�q�5G��Юgm�9����$��55��ݕ��Mu~���	U�����f8!�d-Ie��'ރ��T���4`Rw�r86�I
�AD2��!#�M�������/$W�ǒ�T��|�BE|�࢚̚�ך��uF���Č/�!���"F�����p9���z�~�x�J�Z��1(.���:��V�0Ll=OR�f�C�����r'� ;rp����>@"ד]�i#�|�ѱ�[�6Z��P��$�RًfխPh� �EFR� �.f4Q�p��`8�?�`꧱�xX��7][Y�f"Eͷ��V���j�wL}�OM����Rʾ�!ӕ��k`��� ��z�q�	�e���硓�m���}���m�g߰7�>�,J�2��G���8R��3�?>��DQ�e���!ܗ�TL�MO|/{ayh�ҩ[F���XB�S�	w�a7�/�!� L�>6'P=��)�p��O��%!T24��������+�^.�i߀p:.$3A�1�2im]���6�[ �.�55��*�I��^-
FQd��n���ǰ�[�ͤ�Zrex5�����+W�SWj��@ȣ��S�O8�k`���8����)��ɮ����)%Z <�����+d��3�6�
�~��ڄQc����6]ٜ���k�sr��R*A{���G-�,lد�Ajx� |�"�S�T�}m 0���L��n|�I!q�JWk��
"�/��Y��ؾ��
�(���8yH~|��v���v��.�D59�P��/��n������������_td?�"�X��>�*����a��� HD��ޛ@?{-{b����0�ٝc����j�x��8�=��o��1j-o�9 �GW�p����/o��9�#���o�Z��04?��$6��T���
��>���VM��;oO-�C���/�,ŀ�ҼI�e�'���2��K��!��?6��ɩ3<��a
�@���;�K����n'F,��d���#`#[A8;,�>��]�4{$�>\���|�L��.����'9�E�.���R�IQYSE���ą�ˤe��S�5�Kr�x1�2N�S��G�ቫv�\�[�>�_3#��S����%��[(#,?�`��%�\�	%����*�S�b��ZLY�Hu�n�o_���(DyQ�K.���-)����1��$~��`n�U�׋q��7&:�W�ֺ�"ꊒ���� !{������0��^�BU@�~�Yn8y$��Dt���*�5�����>�"�Tʯ����*}R��9�=�I����<`z��V��4so8�D�f)��Ƈ^�\|޶�*̧��,c�- ն�܏1l

S ˇ?\����T��2ƺgu|1r�%g��7��]�Sh�Dç����V�� �FԋNA�^h���B�rs��x�#ol����OY�\�f�ZEfx����~8��W^���	�T��
�bd<�����\4�h��c��:��+��a݃,TNB_���i�V�]�$�2ŉ��ږ�k:Uq�؛C�̢3��Ca����U��!��p���!�~SA2 !z����j�s�D��JLAC���� '�tlU	9�\~}�,R
vEa3��d33TN�ԑ�Mk�21c�I��dV��������9/eP�� �֮�aC!�JOQ����� cT�Ʌ��>(�O�Ь�S\}�[�]����$5��Ӓ^��BA���2G���d2�䏹=��)߸��8oQ��NF���m rfl�g>J�����8s��&95�D��u�z΢�� ��k\�1 V5;����-y`��t����C�]bs��P����$�gV�B���k`DP��O��[��t�c��KGҚ��(ޫgO�sjK^�(���R�� s{73*�MJ�m����mA��_O����`K�f�sa�:�(H���J�=Y�o������iï����w��o���$ Y����(U�{���%8�a���y(�����=1nu�f�� �������A�0�/~/����,������}90���K.�)m�\��nf���{�v��1�:>+�X)���,K$tKvs�!.�pBvj������U{~wkU��!5����Ȑ*s����`֌��cy�H�-�?ç�X؆��Y|��GGK��)k��O���+<�Nr��c����O���[>b����[C5���#��������괤gi+@��-TVs��N!=�<䨟�S�U�t�,]�Pl���6�Ⱦ���VV��
_-�eā2A�&���4��$�x��Փf�9���ӫ�C)#���I~5K4}����|�(	"��V�B�^	9�4�L�B5wp�]�1�� �!C���5��2�::۸�=p������h�<4���uv�If�j����P���j��wۑ3��*�8�Ī{��6Ŵp�AX�J��]K��U��~_��+Sf)4i.O��*d�Z��RL�M�y�h��x�a y�R��p\!IQ�K��k@э�� �u�t��zϜ�]js1p�W)P�ε@�a+t6�%��VD/Z��E�,�� ��b��Q�g�G	�r�.>�w}�%π�#�i��sH�Rr�������<����hx�10c%X�Ov^q�9w���~��gmQ�x��^kg���>�Q���������x�GAI�s�}�����f/èE�P��-���I��~�oJ��#Zs������\���O�N�b�ç̱�2��vh������v����5�0�e��~�5[�+-'�;��^�wV���a���	~9=M�]t��R�֙��(�r�E���V�GЇs��ds\l!���x1Jp��XG2\c�u���Ka��n��K�0?S�f��č���������}�\��qԫ>��M`g�wϡ@c��fwygز�~��!��w�%��!�"�PA-R�BX��:�awҤO������7Q�t����� ��&	�b��^�J��D�����A��L�Ll��y,����`|����4k/J��{�rx3P_�L�1�B�r��K�XO>�un9��� o|ŧģ�1�0*���x�!�5t�qa~�#q����o�������[]?���6R�w�Ѽ
 �����y �P�����0h��)��f��ǏM�����2=o��N!�M ˬ6[l�E~*N(_�C`�^�I#��J����e�th!U�v%�Yơ��ýH�/���u��݆zU K$��݋�)�*-U�RJ)(z:�o�������P���?�� �%9��І�s�t�����o�
$gn�nDr��&�,yD�T�W�]qN�2�F�:U߾	n�����Jb���gxH1�ɀr�K��MC<2��]U�*�E�q�撋R��049���t��UG�C'ۉ�_/o� ��˗��dl�r���M�z�S�=��N`ҦDo��og����!�^i0<l����1�z��I ���K�h��K���i�]������ ��K��`��'w5/�"��U��~���Й�C�)g�}\������D���Qg `��i��)!Pۥ3�N�>�2��9EK�-��g�EOkζʆk%$W0�e�[�$�C�����3~�����/�� ���g�����\V���v���D�!�� ��w����#�SFk[�^���6� >����<i�x���H�7��ve�:R{�	���:�թa���]`�u��%?b�<��q�Z�hER���d��=��r�]a�
@��3}��6�
T������a?���ϮC�4Q_׭��)�ఔQ�D���+*=Τ���^%<yª�p�:ڄ���{�3�U�89ؿZ��T����Ib�T>jpd������S��Z�q���#������=��8��D�i��Z���s|�n�.%{nͯ|$���H�gE�z�6j)��Y(�KiY�⏳E�B��*Xg^�_�)ET0�X����f�v�����J��7n��&��+-���8��t]�ƹ�E�����&�6�����!4�-8�䛥���LDaW��?��AYwq��Ŏi�&��������t��j�J��b���)r|*d�No+Is���;��wO��y�����W�� �D�{l��ay�y;<��[�i�hA�xC�)� ]����	���	P����Q=��r"��ǈ[�ɥ��3�7��5L ƟN�|bq��]V#���Y�A��s]����i0~�'�sV�qƓ#�ko�y-SbJj��E�^}�}��&q�_��M�>V�$���M�ݑ�tA�[�����I=R���<���h�21<�r+�5)��wF�&h�=l�Z|$c��IY������^-�	��Ɔ���_�˓���:��揬�y#<�im ���2����A�).����UK+�c��,�V��qW$����E�o���<��m�+s��E]����������HX���.�\��S:aD	# �A�I����2Q�W�C�i�.�����_t��t�JHsQ(���SX�~��i�N2Q��29�^؃5}|�����k~�3tr% �$�|$�����B����P?3��b"�{���E�?�Dn_���
��t\)�ls�@c�X�=u6��9�/�(���$��ʶ�+��Et̶'?��FJY�m��1�1hv83f ����0&$2}<xN�&+�������Zˈ�_4����̛&��}�;Җĩ����^|���z]B�.�? �k�+�a9F��R�|�Ǽ�Yޡ��T9��=fZ�u�|� �qGn�����2x,tq�"�]����{�Ȼ6Rtjm}_L���v�q�Yn��h�q���g,;�s�g�t!�̴m�����+۔9m�/�e��i��m���1�6�����C��А^��.�p�!��M�l�sB�Ѽ��1z�֔��v8��=K�7��~��..�.��	2 ���h��=�4�6�{�',�x���lK�A��ho�����Q'#��g0���y�vO��.�48蠿�Q��d26�?J�c���p�\��bT{y1}����ʎ�V��ԯ{�]?j#�@yF�m�Ri�8��4:��I�~C����\П���H#p>�Y��{3z���)4b{'��_�L�Rh�mF�/��ng�gw}������A��sv��0�I���H/ Uo3P03j�X�����5
���w'�Yn�X&�遼�O,�GN��Mr)r`%z��ZZ�$�3���V�����|��ey��!X#"�a��P0�|\CzVt�S|u6}ȷD�mo#ʐ���`����lƏv~Q������o�O�6��Wn{����zv$�GG��� �Z�rzE.�+S�
���`uԗyU#0�JG�g�X�/%�И�쬵�bV��[�H*�F� ���bK�X�5/�|��Q]	l�/��B�np@?W�����46H-2l���\
�!�^Z�*�Ἴ�0⋮�V.o�3@A{��ٚ9��Z�#�6#��T�ҧtv�KV�'�~���Y�2���hh�%d�D=�����J�h���j�	*�Q�h��gԁ�|5.�d�-[!�՞vH�� ����e{rn��(�?�c�s7w�L ��z��/@���7�=`��Q>�k
Nl�L���OW0��
�����H��t��J\*��
�Hѣ;]"�P`��if���m���pr��R����,�^��/�+�j[��	�b�#���g�U��CJ�ZhI%����Z��P4��ZZ��z��>HX͘ �.�u �Іl\S��oQj�J����5VkT�:�B��ٺ�n�@�����z�s��|l�;F�Y��@7$̓��La��:ҫ���I�],8�W��&ěѸ�������9�vR.}� ��4���M8Ck �������
� �'c�ʎ�D9��(��!,s�o!�3fڏ�����%㍄r^�sxK�bU��̀�� iGk�K4�荣 ��lxs>G���\�κ����>������ ������le�唙�좭��<�쿤�2�H�Y�O��j����iX��3�K�v%�r?qK�.&L!�/e��g��B]�e��>�DC�x�l�{����\��Z�T�5I�K�U��Q���6HZ� ��v���9---�nqu[��9OV�`.�$(~��LT�{�i�Ƿ=�Ѵ'0��5H�^�b7hQ%�%��/``[7�]d�2��ڕ�w���YW��ry��:f=.3�<�:�7�� 2�..	z3��F7�'����!J��u{T��5��[e�RWvN�T�K�/��\X~��Ah5�m�q%Y� +�
_`�4���=M+_��{�*�y(\A`�&X
�v�~�0�v������y����t�+Jj\���Ww3�dTl[TޯCAo���}��~P/$�Q0�9QI�Y"�5q��11ڠ������K�c}I������1[$�8����V�]�j�ۿ��2��e�RA|�����]:�C�TO�1��]w�K�1j�Lpߗ���9@� �bm	�� dy��aU�|΀��6E�S!P��"�	m�o��>%
4�@�A�N��`w*�#.��Ea���F�����C���')\���X�~˙܈�vJ~�4�ۣn�!�9
�_^�Si�!n���$h_	���浮NG�5���X��u���_��s�ǐ�1��tQ��
V5����#[b��m�j�{��"^�U(�f2��7^a�/pj�_��o},.�1�&6���ζ M�C|�`��Hү�)�KD�3%�H��q�".���ϔS&<���8p���a GJcn&�tg�SC�Dh����K�<!��L).6�	��f#Nz@`�{��<�Vz�0d^X�*�?��Z�$��u�u�k�E��P7��>!ܻ��Iw��X ��'KH�&W6�f��
O�?�g�5l�%Q
,^��})N��@�cA�;�1N�U�ҫ�l�Y��;�~}�&&Y:R���
��hck��2�oz��q]%p�i{�FK�<�1�P�Qyы <���X�cH���W�A�����gکYY;Ǚ�Y��huC�u|�_���ؖ�4ħ`�Ky����Xm9�Yi�:�T�1'��_��c�mD@��DCr\֘&�J㘀縜& �:�R��Ô̲�,D�{���%WC<�C��ku���K砠ދ�5?N�3���D��y�#��Ǜ�N;���ܗ?ߌ���<\������]����m�`��a%�k�M���,ZU8��?��!*On� �GϓQkR�����x5aNˢ�G�c��dg�z������#�����yҗ�]�c	w��y��ĉ������&�k&�u��<c�b���L�y�%:��U��@{c����O��5�G���_g���|l�p7��3K��yE��4� ��U�W��V�O�v�K�z�<*#�A
�N+>"�wG�y�Rx�?�.�i. �"�=r��F����ڮ�I.	�M"Ql2������"��]�nhy_���<"������R4KʝE%J��O�4&5��=�6;7F���}�L�;���ȑ�� ^�H�"u��������������\��U|�I�7܏�k�mW��qC��]z�`2��/��#v|3]��F8�^:63R�Ct�pə����Gd��h]�:�*��g�,+�}�GӁ15��ѓ䈟d�ΠI��"�/\�ԅ.`%����>I->1�n�8����)�Ȫ1GM/}`�$�n�,�� ]MG��_����J6��^��b"��3vշ�Y��l����Yo���؜E /�U��%�Qŭ �"y�7kt]��#:lIq��-�ym��ǌ�I�K��m���u֓�SBq�m/�'7���L �h�Qs:�B�{u���ē-�G�A,��p�mUD�"E�=����bq?��ak� |��D��LԚ˪&c]D���GAC���S$�`KO�=�����qaH���Ͷ�Yo��-����ض_˥�X�i*���"o���s˨����gɚ�ó=ft-;������U �j�t͵1*������,tZhR�w ���{h?��5I��:���U6Y��[�kn�4
��j��h����9M'NL^ιN��!����l�ۄ�9��v(�a{[��۷S���E ��Մ���D:O+å����=�jW�`t���pt��|���C7��Y��f�2ѵ�8G5�hʎ��cF/A^�:V{M$?ݰ,%j;�m�E7Ɍv��М #��>C��ٱ��Z7�^i��ϖ��=H4b^��i��0{V<B/�4�2��c�zd�Mad��2�I���̫z�rܗ��H�C�ڟ��	�}���q>��Ь��A0�0��)��[EhE���XL�6��ݸ�x�����T�sitd�l/a��4!9�F�Q��?�eU������Z�<�>���Q�ڶ#�+#��_"L��DU�~̗,��(\x�>h
���0pcf��HVҡ/C�i?�fnU����vw�ý��(�|;�h$e8�����$�<�r�szga��o1vǚ0�V�j���pg�5"ս$84�ʏ��^�)�R�1	+���n����	�B�is6`勆d:F9�;o1۶b5γ�r	䟣$���C��@���gD&�:"����,ӻ>&�]n!ux5T+��RU�7�A-d��@�x�U�?R��d�v��=ʨ.m/���pjl��l���WI֐Ü�]܉�v������A[i��O،�7I�>�����4�w�b+{�ȋ׆�@{���k����&;��uD^����������K�>��B�n�v:���}!�:��~��Q��"�NZ�{�TQ�'T��"�&7� ���ܘ�a���f��2a�I�>@��]�e�H}竰SiIg���m׈����USD�g ��sX����Z��F�Kl�Z�QO�ι=��
m �R�H������F�g��[�r|����3od��HO
��5�D3�ož@=^H��s��~'�W��b=���m�h�������m�@W}R��]x��1A��������� o6�Sܐ;�pIOH��J��		t����k�G(L���RA�y��������"����R�����S�K�Y��CPYLy��;����(إ���֙e�#{=����>1���'�_�v?����e�AǢ��Y~�rK�&�����\��̀MM���Fg2�4������%n�i}ǃڕ��S�ɤ���NvR� b�H�q��c�e�`�(�������f���Ż����p��J�(���I:�P`��B�O�
�/E�*w�o��W�Ѳ%[u���"�)ŗSl�j��P��f�J_�X�� 0&��.,~ں�WټI���UƮ~�h�����Z�_�x3����P�n8��?�����i��=l-�F��d���ȶ�v�c�`/6�0E���xZDj�*��p�$�\fT�oy ���l��,�;
�@G�XN���R�h�P�9�7hBc�AhG��9'X�	��䐾*!r#�c���B8S�Y �{�ް�.�r��R^2�.�x6�)ӷ�9��Fz|!����i��n�Rs��_�V ����i}]�c��R*wö*�+�n�:FB�u{�w��;�BY"9��6�DV;��_ȮV�y�����&Iǭ�M����U4P��,�iȹNSs�[��No_��!���`�_�t���}*�����FΉ�
^o�[g�gH�di��~�%� v�,U�(��m��mj9��PVfg�%?L��Y���3�S.���'�4�C���d�Q�o��qxE-�*ئ���kZ����d�v)���OV�G[Jysk�A���Mmv�Pʌ$�q�1��e��&�\뢕-C��6��2x�Y�QC��|ދ�k�"׉��"���g�����K��D/���C�HW)壘�����<��g@�p�5G
B�{��h�s�H�����#��	Ow����ۘ��'�I��6�|2�f1[QV@�BL��{le�BB䗂`1��6Kv�G���=k<�l�n��{,+w�}ẍ́Ճ�NؔOEY;N��K������ 8�������[��p��[�]Rt΍;E�K����)������<������jDG_.�o��&�u������� F:th�Hr82;�.}�{}�o�~T� 5�{}9�$V�E�G$���Bo��G���?��U�;G$e�ԋy�:Vl����^���4H���I��Q��1l�`�r/�`�Lp|c)�yN��Ԯ]ew�yFaM�%�ԃ�Nl��t3t�>�1� :&���o���G���Rx���/N�>��1˂�1f(���#�{�H(`�S��)��dY��>X�7����5/xʰ�� ?�b<@{�&�a�$5{3�?W$����f�l��;��A�D��|��-(�@A�vv�ܠ� b����'҄�f�d�&�u�\������GgC�u���x��Ŗ�lxcR��.E��h
KI{O^y��I�8��ũ�ci��_'��6T��wQ���i�*=[wk�5���s�"���n͗R�6��U�KyH_��Wц2����:u����d��w#���/{y0n^bu�4��$c�¿]G��9�7'�J�Z.��(�ԡF��\9��c�/xx��βbC�K�p����;A/A�m���1X� �+��[Or6M�$�;�6Bx`�|0��+�xk"�g$G��L\�ZC�27w��[�/�ñ�C��CW��&8x1��:�@|��"��|����½��q'�$���a�7rs�V���J7��gk��U�V�RƋ[��6	��Q����f�iº}ժ,�.kż8�9D��SK��7�Vy����1�%�ں������B:� ~c����I��G��~��If��:�cp�G ���o����Q	���LZ���\3I#�[{�;�r��#M����/��Cү:����Դr��z�P�)��1jAgp3RA�Y�u�����v�w�m9 �3��t��ߒ�����ډp<��c�o]V�vTu��ax�j� � �u� ����*�O�$g�pŴ-Y�s�jK�k��
f$H"���/��~�\f k0�b��GM����=�(m�`>���(,� �E�����z��W�|D�	���Q'��.*Y&8g�U�i_�������v���( 8�]-
]�c�&����o�<�J��4n�)��؟h>��'��M]%~?v�C��Q�\X>ϫ�1�;v~¢Qcrr�����@�O�C@�wr�6�̝�-c}I���rc�dם�g��i�a���/{M��#D���p1�נ��)�s��4�	3�E���of@�48�G��#���9̤��L^L��vb*xحs�k�X@��#�u�euv�S��V߸��U���tx����\[�N�!M�����_}�����'�HL���D k@�V��'��g�?�����6��i.��P�?�Bm+�d 
��9qD�D�B(����{'��(��i�R)�A>�u��g���ӗ;���>�x	n�du�g�Qs�m���d��gG;4�@�:W�Z���=�������k�L�*Ej�|���|O����ZSm?�2��������]P�����/_��-~��Q�[�bdF8K�ϊ]ӝ+�*��n��[#�&vX�r�4�f��]��pK���[��@��2A[�&����m�ћ��7y�q��[LFka	�Nx1'tu3��)9��Tg�$*�'uez�t/���vi�@I�� o��E��iҌ��bq�k�>�+���I�0���횏�%'�R�ټCB��ک�#~ۚ�PbxK#>����O���=�����FQ�P��h
-�J�RxAG��I����ٚ�v=�kӛ���l�\m@��woY����˓�5��@l/Lh�֎.\�y�]��g̗���L�T��IP�%�-G���Q����(k�r��J<%���5"�����n�r"R�Y���#����ؿ�=�ܡ���!�x���D��Wh���D�̃�CW!9I��L�U�}')�Ē�!h��j<<����ڕs�me��B�Vg��
ҴlR�����A��<;ĶV5+h��x*(�]2V��eS�z�Z�0�H�d�����Zr��spX.�hǫ��J�q"��2 roh���h3�@���]�/�d�~ѵY[��#����h�d#�$���q9$��#��P*C���dG�H�}B��؛3�EP�O�0�_l�\	g��K��O�����͎�:��-�0�;��C����K&��jAw���Ӏ+_���&Юh��׹���%6#���둞.{(�7��-�1���ң�)I����1�U`$}���a�"�Qs��K%� \2�����1"���G4��[5��I���7����F�sV��ȭkj1�@�+�hG/{s׋a�F�u&iy�5 ؛���0 B�6)�s� �6��$`�%�	>�J?+ ���i�����MP=y�N�ѾN�s:�%3-IJP�#)�JڙP�%�Bș�elI�7�$�?%~���ȅB:�y�Pl3���e�1n)��^�3��2�*�!;����Iv#���Ș^����0�ȱ��کf1�?;ɬ�lR�&�Kp�T���`�E��N�)'�?�<+
t)��|�Cy{�0�f�o�Ci^;T��CX�A�X1�d�ô��7ڄ�j�G�Z�vG�o��=ӠL]�R��F�VmK��+;�؉�zh���F.;���]]6B-EF��������N���&-�R�i��
���.�>T�R�sl���Ƌ��\��}f4@]j �h�ߙ�#��g*�uR�V.�����%Z?]�>"I�%�T p�s���Rt�U�{����A�OoEG۰�ϝ��8����o�Q��ǸL�<�얨���0���⢋l��^r9#�vGHf ����
��Ȍ�I�D��c�z��=��D�)m��FX�3�0�$�!���\b6w�)�����X��.�\f��u�2+�����[:X�b ?��~�_��UQ�k��:߃���k`�wC��mT�Į�{}�j��J@���~�[��z�䔲��i�,�v0ޅ��'�O�ؾ��=^�'��e)A�Յs���ns�@��¸�gb���n����V�Z�
X��\��t�.����(����\��&L��?r��� �-�v�*��gu rH�|B��ġ�~�<��	��p������-
��D��w�$��g����s�M�����	qv��8��.���3��%њi��u
�L!�+(S4KA�3��ҚW��]!�r��cډ|��-�æ���bJ(˔3�6=��ٟN�="��&�������P1FO�ɶ�������I5#7�����8�(�����+�>�7�T*d�#��܊�Cd11�ϧ F�Y�;	�K�!C{ yvgm�'��?��)R��0�ZHe�,�⹅ES�w�A}&b��Y�e�ة�BN�/�n���tgJ.}�$>�]�4�`d�[�@� ��ÇI��������-��7�!�P1wc)L�C�H��*����!	2�;�p\�R9��=����m` p3m2$�h�wY��>i��ui�8��s۪��M��*�y�qK������9f,�5�a����/ 9����a���h`߀��0O�ja�~����ل�z+�+��>h����~��l�~AI#���f����.�7���j��#���Q�ʤ���%�<ǰi3��CiȮE83RIb�ȓ�a5+���!��N%�������ײ�
?�;��	�\�e0�0�f<v]E�纲&e<�c��z�M��q�T��CУl��/�h��pY�XY�u)s���x)dw�������H��i<��Mub�nhl
k�0��!w�(2����*4����I�V��X�)=-!	����F�`�b"����-�h��w�)�+I�bA��js��
��ѽ�B��]��;�����)�i�p���=�UM�EZܩ�j�U�:�zN�4�\�&
�Sz�%��X�Br���0O��,TC�
%�\�E��^lf�3�e^���7��
#�4د����&�k]y�a �	X0t)d�]������-����!����]I�O`z����};��W�uX�gV�4~������)�3nct���s.�t2+��@.��.���m�U���=��t��Hʊ�o�X�h�QV�k}������w�L�AmJ��С	^(��)��xi�(��� Ja��OGo�'�ĴM_�G;I_3IY�����E}���mzx�i`�>u����d���l�m��a!�6H]�5^�0H]�)�qG�bcxo�A?|����Q���WlF"�|=�戴���zˏ6V�M�w5�]�Uu[l.Zh�G��u9ȵk6����Y���E���l%OGe�x�1�B#q��'Yϰ����!��wKœ{G���>������K�U��M�<H�ɜ�p�_��
�u�.'���L.�)X�c��>�wlP< �w'�nϮ��+|B��7|�~��:�_M�͐ɽ�5�9�xˇ��r7�^����7���g���c����6�zG�T��78y�+���t�z\D��AT�cߴ����6��4R_�<WS��4����*�\Ģ&&@ .��򜪿Ǽ{�|-��C�`t�Y���a�5�q���-�i�O���=@U��&,�&1(�����P���{�l'7ZsV����w�D��l.��,�z+�K�TC��c)[�� wBa�����2l���3f�x�ޘr5ImY��k�����Uq���Wi������I{<�v�?��x�fY܂��.�9S:��d�I$�G�fűٸЬH-��jF8��7O/��ea�3�d�g�T�����E�y�O�9�b&`���Y���X�]~���,&{��l��}y �J3�
�C��-T��6Zr<�*y[1�݂x�ЋP_�	''RJ���Y +��Ӧ�7�j��Ci�y�71�o��L�H�r���4�6������c�4���	�ڳ<��&�(hQB9����^��Q��L�R�DV@-�ܠ!g:<�\E,����n��P
�u����S����z]�V��>$��x�{�B�I�9|�=��6	c�� ����&��J�7G�L�/v!l�bhWX���{�K�P�e�������z�+Z$�sj�]��G�;��Q>٥MЯ��]��2'�!�xJ�6Ci�/o"
�mk��G�O��^�ɰ$u7���$��(&����4����U�����^w��-( ͤ���VH����. ��oV�y��1B�~�@�~�C��V%ғ��W��y�ƕ�tYPct"�Hi�g0;V�,yYu7{J�;̗�Q#}X�-��)7T������J�k�����0G�ʤ����¨��Ȭ,T�����7>����N�׳-q�������Xe�c���`��[瑣�BT�Ж�Rv�%��T�"�Ƌ/V�u�T4?�R}q�b3��}�q�P��z��zo¶���[�g�,�f�'M��vچ/�\p�ܶ:�6~_�|��+�o�����
Y�e՗O{à�{ �7�����辮�"���?�Z�w ��!G�^5�P�]'��.�&]�B�Y5Ȉ�̬��k��pQ���ϐ�n�+���\Y9k��)����\g�l)��8���gO���c�����/��arL������6�Z�?�i��Ә��mGX���`�w�$�h��,���oԎ�7R�x��ط+�C0��]*�F@i��	N��LPz�f��<Y�σ*���c�5�R��vP#ݖ��G�K��yq큩	`�V��˭u�G-���5^���[�ݞZq'�b]B��Ɋ��:
S����T�V�`=^�x�Ӱ�)�po,�Uq�t�M��6���1�'��R</ܵH���V��1V_�%�w{���^�T!��!�>x��S�xS���G���{f�w9�<�Vԡ�
�y�nވ��{*ϧ����RuJ#J�ܽ���M/c;���?3��{,�aI�#�g��,?-�ֲ��Oҁw��*�(�=�����w��:Hȹ��K��CqR �`/�7��^��m4S�+��Fwɏm�m��H����l�m�R!�E!Bh�ڲ�-ͦ��?\�a
�ϰG��_I�pqq�}j��~Y�ڦ�^G0��q1w��`�Uv6��?��Ûd!V���\�I�� D��� ;�pFw��k����;'�tQV�)�⮎��*�S�bn'S{.M�`e�b��,��5�����n��2.���c�V�m_(-���ˀ���1�4�6轨w��i5e����JF�}n�~va���>�%����c��e�Y�su"�*G~�q\`M�viŭX��O?B�H̘U��M�$�����C�����R��s��T���Q�L���}���x��骜���K}ܨClt�e��c+��cj����^���@q��2=OD'�l���C���!`Kp[�	�+��Y�0U�8'�PJ�~�bQa�@�^�v+~ϡ����5��4f��[��{�����'Uyl�D�s�h^2�Hd:�];z��XR����4�+,i*؇g+��,M����.��_b���-ϑ2c ���Lw�fr�<�Ǥ���������Uш��I��)$Q�f��R��ĺ�%v_E&''�$��[W,%��G��1��!	 �73^l�鶙�O�m���a�B)����{B����	��/&�Z��^����nk@4�dO@��s�v"F4���5��ÒtEg����rȸʺ�n�������߫o��xI?�zZ�$L5hzӲ�4m��Ȑd	�%���	/�z�o����o���YB%�	!����OΓ\��\:���g��h9�d���me�@N�E�y]����b�8C��:�nK�Ls��<o0�����^䌞m��#41���;42Q�74Z���*%��)|��پ��]q�&��"g"CyΊ��'���u�C��z>����v�Qy�)^R7lJ�<�_���dNR��G�,r���
��}�k�0�\x�%؁����������u�\kֻ��2��-�<��0W��|�N��g���?���y�E��3��l�[��(U0�C�B'�%aS�aFGաxO�6e��>�����u���h(�N�Mv`Efp.�]6�H��Q�h9����k���^��U}�aA�{���Z\�D�{,ishzU)������:�Wm�k]z�Ҥ=N�o�X��<��t��p �-�n,r�������l�]�������H��Q����7��Yc�y3��=U��ξp�U[ٜ�c��JKY�1���LJ������1���Q�m�n�a�X�@2��1���v1&N�R���%�e�FQ/���(�~��)R]���^��vp�)1��ū7g�!ܔ}3u��>��e���U^� Ԉ*���JG��c� ѣ�h��%�d
<5��'3�$�<���+�;��5�j3�[�a���gp2/��C{�A)�7�N���<S邑�FpqO乙��8� � '�[ !I �HPcBC�L�^|{\n���T�����=��&��<�*1$�̂���xR�u�"P�}X��a���E~ES���7+��p��_\Vɽh�%��.�
�u�e��$13��(����x��$a?�JU|��O	\�t�gW��|�}ڬ�;R���'� ��4�/��C�w�`h�Ip����*fJaK:U,g�����0z���ʙ����2*�e��>B�u�[�"�Ř�ʘ����?�a�s���$6-�GdH;��@�[��C�y��@ ��"aD� !%��*�eRma>�VV>%QX�Tf����P�k��?�".t���1sX��V0��ڼ�~D�2t��5��GQ���{y�v�S=��hfC�٠̜+jdpL���eS�|&zj�l���Ċteр�ʃ�Ǟ�����/|��3*X�
�[�*����1��$!���2�LԌ,;4>Ť���U���tѶ��XS|�N����i�0�3ׯ�h!�ň�p՗�7
\����Mk����>�e�P����c�󁸣RGn�rU{#ěv���r<ʇ�	�<���|��~���Sk��/lx�Yf-^��kW�k�W.�$��@�/��D��DL]YgG��qkq���_��c�8�̽I�b)l�ܔe������mɘ��qy,Nî_��0sUt>t�T8�̻/�!���e�����L��>X�2�s^b�a��@����}~tE�ן�ko���Ġ8aOgNPR�+�%?���*��o�t6��II\k�ň�i.'��\\y9�	�3�B���|ЇLl�]�Jv�]�ȩ�^)�a�%�r�B���(3��c�G�meG ��@�S����<��t���E�[�0���2�O!���q����r��2�� �&:���f��|�Sj���D�G�_��C����A�4�#K���x`����l��>ے��ے�����A�(y��mD�+l��Rp0|�X�Nm/�N,5�$[[��a��W[2�6C Jj��Lӛ!Я=�(F��y�mq�� &�2 �c1�MmK�[p���v���SK}�=+�e��c��bh�UZM���"���9^��h�}���~ʙ��l8*Y�1.±{ �F�g7��fݤݡ)A�P�͚q*���p�w��T�{�?a�����ɼRάz9m����l;7��]�t��R�6L(���ٷ&�A�Dn���t�v-\-�_�z�1�*O"�Nv�;c��2�.�E�0MG��jz�� +WB����Tl�����v�C�x�`*[t�]�9��{��E�Dl�����p=j�5-X4�9,ڮȧ���Z��iki�+(�<Iɋf��F�$��j"�2h�)Dm�Jm������g:����ܩ}EO�Ls`%#!�s�!-5
��B���_C�:Y%'l�`?�v��nS%v����6�0�o��I�qJ��=��I�0�
���H�G��T��(2�3�ئ��:)�p�2��T_V��ǖ���}�����|�@�'G�-�-!��:Q���PG��:�Hr��C#��zo�Z
���,���{������870���o�ȐF��"�d�Ɉ7�@��=�w� 2:@��+�U/ӫ�Y��xjϽVh؇�������S����9���N5/��!�+%��[�D���m.�W�Kf�8�[�L<4�m��.k�c��*0�'<\ዛ�� ���뽵Ϸ\�_G_��V���	��n_�)��J��	Y.�E��s[��B|*Eb{�{"�F���]�0�~��v01�GP�4�[V�Hn	���)�U�*��ڷ4}��Y<x��a�`Ю���� ��8�|�V��u�����<ƣ�*p3���Ib#_�:�����Gr(����mӾ[=����}�m���'C(��*���Ƭ�(_YC(��/���bZ)M���o��Jy�;�nPz.�ȈX6�!#wK��̾�˺4o��ݎL��p ����R6HC�J^����#�s�8���k���~ɇjo{����ng<� ��Q_t�5ش����^H�$	v}Ĝ]_�t��&����]G�x��WZ�t�۪��X���s4��)d�$?������X�S
�+�8ni\u�aQ�X"� ��E#K����S�G�a�H���s��=2j�qsb'+o���ݝ�Ϣ�pmf
�L��O�D���N\���-��y5��$��2�����t5}��b����PzA�Z������m9�V~�	1���XbG�kύ�X[E�%qW9K.|K��� B2����F}�,t-W���R
u-A��{�����
=pA����p��V�V��R��M�ȗ �1��z�Уg!K��t
�ja�f�!Pv����T��&�`�1�ʄf��ƙX�_�f,�̵���.-�M��'�q�v�Z��Bg3�_��v����} �U�b�2*������HA����FO���IxE�\�r���P�X�&�Ϫ��rנ�>�7(
�G(�˳��h	�"�fj��>2yS�^���l�2N��	B��{i�ʥUC�7m���ÐC����� ��{�8S��i�*c�0�S&�ɷD��ר�4��������~��ir!z�6z'Y=b3j�k&.���"�h��&j`��DyN'4vx��_��oE�4WF�"p������L+vA��>�Ӗ;#���t�x��j�5;}�.x����*%�Ԭ��~�!3�����rR�L�a�jWS���+6�����w�Vy;����#~7���n�CA���{�'����N^p��φ'ik\���O��Y,G�$��z��!4-j���0�=w����d����0��9Y�P	U��1Ԛ�����oa.%���T�je���!�8��,y����Yrjò@���<�o\e1T8�st��"?�,0ĭP�N��H<�� cﳓ�N��\H��Po�lɩh���H��� B�1bw�j�AI��S )�6}V�4?�a�]�*>�� �A%+���>������fk�?F��������'��BЙ���Yy�*:6�[f�����XR+DH�_��B}!�[�{�c2KS�Y,/�*�^{�6�N��׸� ��� G%��[0�jf�S)�� �?�J��lCsu��z����=zd�J���A�=��$�e]��Q|zCVX�p 4Ez�R�Z=���މձ��ba��*���HQ��N�5pzܻ'`q�	���+�N��O:A<Iv Al�;AIY)����?dv]%����wU�=Fl��!=���R� �$� 姎��Q�(QA3�wd�(e҉�%Y�5�P4���]�xS�����ޯ�ɉ�)1ٳ��q�aР�
�+��9�T������MV�e����3�7�z�4p���<_)���+�����c�=bA�#�o�X7�G�%O�5�Ћv�;o�u�Ֆ^����k�˔����r��R���l}Q�g�� ��^**��+7�깪ćA&�!�J�8�,�{@{��󣜰�N�Eh�V�g��c>^��_V�#�rv�C�#Ƭm̫�5i�T����`�f}�Ё�~E\AT�� �� �A��-G�e˱��W/�,��=��@Sэ��8��'}���=偾�T�j��F��I�*e|��䋳��8������3��������ۿP��š�q��XR)K�������(
����6	_�g�����
x4����Q���s+2"���`�e�y�c��upˉP�盰�gb�W#M���J��sJfwe_
�����I�48����~VPPj��<�����~�#�)�<b3q�T4��aU{Y��v��L�'�Y���|bA�o�c�X�#��� ĕ����UwԄ���X#����`1�v��.�#�T��@��N�ɞMܞ��x�i���*�@,*Y^�|Y�&O�@���p��;���?�E����@T�p�6��j�0�mR�Kw/A���$��9
�����%�X�c��H��̽�	���������Tt����9�6 c`������Pؼ��+3B@{[���|�BŶ��%���7�L���(�^���I��5�{�F,U���Q�k:��s �zw����o�y�(m�aj0���1�m)��x�q[#T��ԕ@^���Mg\��ʚb�u<#�09�\ލM�R�\R1�0x�:G�sK[���U��:���������,����~��`
v���QA��g�����]>�a�_68����5RO�1��x����^��k�0)AE�^��ȝ| ���m�u��:? ���GZ8�!��x��Q��� o����d�3S9$O[���;Vz\�^���[rS7Hl=lk��1��g�=k0񓁶/Ϟ��CvV��LEm�1@�������u�~T�i �҅�R���������K�Mm�_S�{ ᒐ�����S�X-�ح�*�+IJ5ԁ~���rI8IK�S
���pΦ�]�
v����������Sė5Tk����u���J���^�i�[����L�az���Zmh���׵��b��ק��k�mu���j�ƤD&X��5�qu���b!����9lSScr"z���������,�㡝Zz��>�X�re�Fm�5ӕ g��h������BP���V�]�'���I�v#E6�O_����DO�.BzZ}�cH=�R��ҾG"|h����$:l��X1�!�b��Rir�w�(�����+}3-���O��:�W*������ۆ�AQ��<�ZX�P���VlA\�zIiJ��Er&��gN�g����v�l��?�s4^M��.���0����<+�c'5�Ŵ�z₳K����b�����e6�(�Z�\�F��"�ST�Q���f���b=.��cj7>
�1�U�G���6�篲�Q�r,Ӎ�cm
�r;�:h7Vy5��HՈ�lc)��*�q X�g`�R�8)�Hş'�VR�{5zCX�y5��G	h6=��/�p/g;�iƿ/j�J2Yr�:�3V�ށ���.p��6�����l0)�p�D䢙8�n7��� a�(0�Yv1HiF�����{&%�jC%���A"'^Zp9{���Y����'�����B���&�[��� �\��	j���� ��u�d79���E�Wd�w�"G%����U0!:� U������J�C�����U��ޠ`|W��,�a+��&�T)��?���;�E��[=|��G���L� ��[`�	�ͥ��;t�(U���{Qp�]����\����BvrQ���)��E���N�p�Dg-�������"r����~�3s<��,��%�b*�������b��4�@�u,�zw�|{2(:�:�a��;�@T�
+}�3�$��F2���F�<U�d)9��)`'�-�2��t�	S��8L��7�7��w98͸�}�s>Q�?c�\�6�-�ܸ���V���B�o���-<�
��Ū� cF<���F;`݃�D*��HB!�	0&ѹ���	~o��p���Mn�h�P��x:.@�2�w�F�-������b�����l�z ��W��X�t<P���чi0w��E2�2�r�g�T���)�'���6�!!���/ݒ�^1zƑ���Q��LS�t�m{��N�i���Q�����ѭi��E����9��6�('�1uK�̔# �ejfYy��b���%�V�\����͜N|���Cl�%)B��e�z�)v#M�Usyڗ`N -�wб�`�527���`jjΚ�����;����)�i`hI/Pw(�2��"��4���f�Na2��R"R�0Rp�*�+�4�gG��~,�}r���ib����w7���B�[u/�0{�j5�U, 悦��c���1�:e@T�8�ų��ڐrڷ#*�����ۃ��s��	4�5��l��滮� R�� ���ɗQQ�Э���WU�qF,�!�q�ڼ� .�mg�\{�#�$O-���^6���$�8�Fk�ۼە�wH�j�{�g)1����`�5��B�c��3%���pYu���M�h�y(�����i1�Ƚ���t�@jq�r�箯ɵ��9Z���F��,M]���,r��Ŗ�$^T�)�*z"�\t�B̝�s�ӑf�a�YfC ������'+&ji����Q��-Q
�i�� *�@��6�b��)8�#TO�.T@I=`1���ΜOG籺������K�I AԾ
5o$\�T����2�kW㉡1i5��]g���[�Ihy�o-�΀��O��dZgԦ�������j����e�;*C�F��6(�??]�6E���*A��[�� T��d�œ�3�DK�h�����-%r��~ȑk�Z�!�7��Bv��NO�M�������}Z� %R�P���$���^b�/���P�&?ep9d�3b�Ê$:�����<P.�k�;�h�Z��(�]a���ZC��@X��1�5;RN�:7�ZO���o8W{��J�uV�)C�Ꝫ�#��2\���W�3h��6&�m�;�8ӎ�J�~<�|�������80��а^��ڵiQ_�F�?��M?4�'.2�v�G�q ����P\�	M�^�*��0�i5�CH�A9�����-���[�k��n�B��c���F���_6P���T����U�;��Z��_�P��1�{��>�N�T=yj��%;�-����0Jsکxn���N%j���нB�wN$��?DN�U~�1�Q�l��h��=Savtu�k 	�x=+��׌��Gϭ0%G�q�/0k�����]�8������n�y� eֱ�J�N��r��w���_��T��:���MU�>?�n?�L9d>&�����0&g���]��
?��ۿh"�Fq@yEů�1F|Q�
���W٘Y<����4FĬ��8_��{��8����/�Z�\.�)@���(J��z
N?�g��ss���.-&�ة1f�A���]���yI��AI�]{A���ӗ>�>_v�oG��}A�� ��	�;���Jdh�,�8�f>0��"��j3��Ź�9�2\aQ�-_�QR��.u�:�s�ʳ�W�КZ:��\�$���F][�����X��D-���7A/����3��1��ݔ���b��)%���DǴ��{��ݦ�+�y��r
�kνnJK�a6�MX��uf�=���)#u-���z>[�'LL҇��=�-�Y�aO��dy<�Ȣs} X��+NM�u�z�	τ��
i����f����Q�ｾ/"i4��<���Xr�Lt��Gq�c^7�j/8���Ka'�a���gKf�Y+}�L;u;��m���d�A�L�,�7�P"��]=:;/d��Ҳ"�8Qy��I\��ԌO��~��8����?�&��=��>i�yL.��
տ�"$]q DD�`(?8���b|˩�h���3}c��YG*��"����`��u��8W;�O0C'����8�#�n���V����3ȃL��%�?g�����Vc�wDb`�+	�R�\�8�l^ea�MT����(���Y�vT � PXNB���9��?4��=�����c�h����|�Q�����.��<Z@3�at�I�U�ߋ���p���`�e������S��h�����c�B��lX��)$�_Wl�/���PMZ��
^��@͍4B6��M�fxc��L�^��!�S�#��O ���u}��gL��2�<��[H0�Y� ��2HX��6��R	C��Ҷ�IS$��.�R��OeO��1[&Q�[�nkUp�W�-׻޶��j�/�No����{�m7Vt�3�3�T&�9���F��rW��YQIK&[��oR��L��Q��|�w6k�����$��3�� W�j��0A��H��uqo��E�����v�)%	L�{�N_��z_ $��<&���
}���<�Tp]�}�2z���5��e� ���Y�j�K���n�0�������n`�p~Lv�2J�k�T�+��:颬Vy�T��u'� �ڧ��IDF��Z�DHƋb��ސ�?�F�B����HJ��Yǹ�p��=��&��[݃<�*��W$[�q;��t��Y�&4����司�J������6�e�nC��[��ny�E�>P���(�Y��(>J�U<����A���bqE�Eq窲#q������:S��F��t��^%I�ڄ����h8���.�?��Րvb�-0�Ӫ|JH'�H8'�)T�x+9�O��0��F��f���$oB�Q$����Qj�U=Z���;��{ s���Z��T���U�H���(3����X�����V�\6�׀N�\�=�"�2�x󀚎AƩ^?�م��n�J��e05�}d[p��g�����IƆ�)�e���z��qş��]�X�9�Z��j�]�-���!�L���x�q��7�х�0j���|��g@�L8e˜�Ws�p�nH�A/�yue(O,�
V���^�����8A��P$=n��1!�x�Ӎ�A����*�}��>�}�����`
,j��d�F�2����ivnU����������P�3�ͤ�(1,�oV�U���G�-��E͜~�����0�_K\&)�#îu�_Q:(D��x�Ȳ|��ܗf�g�&=�/0ƽY��5� �.V�:�w��U^x���5lP�ʟSz?>��`2i.�I<z�|75f�\������H�0G�2{2�
~H`Y�/j�P��G0L���tdq����VT2�m�b�\�炤�.��kNxLs�����$E�5��P|(�w)5y#�:e�����?��O���Q����@�O7��4�;��M�#�Xr�t�)67=vt����t����s6dE$��t��@�%��^u��9��yGm����zO��Ȝa�����֕��Ҁ�a��8>- �=�׻��-��4�'��zK�o� Vs	�T�"{ؘ�����]Xe[hbw��`Gou�䚁U����|�*�8TȀv�o�}�o6-a�i�h���Һ5�*0ޏ&'^�V*^�ʕyʅ耭.KBC&�;lw*�.j��ORﰻb���1��{�uzh+�9�s?L��A[2g��9��B�8-c�����)?ņO�YԎ֢�p�����-2��Gl��X�V(~�C��8w<�]Ƈk},{�As��u��ʲ��}��'�nvT�o򰁡FacW\���4m�#��f��O�;7MU�S��;�G��`����>����D�fWowH�$���pQ����_ �^���5ĞF�m����n�%��=�`O�}��x��Ь�w@�'����~0���L�$1A��n9ˡ�f+�c�44�.���UHm�y�D�ҹ1�܍z	q�Y4��;
��-]0D�N�XW&B�4�\OEw�ւ�����	���E�@�HwGA|K�WN[�xp N�ӏ�:�/��-l�YL���:�tʄX�.�*��i��oï@̊
]�A�����f������0�Fݳ���d�I<��@�^��8rbB�]��tcP��_�{M�� �;�
,������KW
XHtW���ttj��B�CZ��'4c���~^ߠ�m^匉88�
�ϼ�(����&�)2�c&A����O�%|�;��QOb���1e�E�wC�?L��{�y����ȧɭ{�xp� ̀Ŗ=�z�|W�����n@��V�1��[��XR�Q�݁�<&�{E�}U����&���aV��tW�;�.�%��
��tf�^ ��x�C M�:rzm.9O��r��l![p���GG�(�qbV6��Vs韡�J�s��>�����tP)�J��g658��:0BP�d���t�]Q��2���Ba���x���A�\���q}�oNY��B�m���,�7_�JzH͑������G�?#��Y؃"'���	�sjG/Z;eE����Yp�ɹz�Y	���ɥ)�3����:����c�����3�uoݞ�(_�V�LSp���:k��B$<�n8�b�LZ�L��?��O�����#5<�ik����rxaG����{���yĥC`�d��%q8��*�� �.-����w��S�H�SW�{&�4@R3C�[QK�rS��꨿4s�J��͓������5�W%1�u˪ fZ��䰽� �PbВ�hW(��=V[�կv٦������� ��"�&�4��ϿLbw�G�0�㊢P���]M�v�`�h3�L�FZ���dN�t���E�UW~���}t�JxJ�w=|��j���q� йx��M�*>-���?J)��0�y��'i�2�ݖ��Cpו,Z.�zF�� ǽ��̄o�W�J4��kMH倿&�����oytoV��g<Iߏ��j������pf�ټx��*���-��(df�qP�y:��8�m}2�O�D���p��:�\*���s�GjY#pu?Z�+�p���d7� l+�r�S�k��L60�3@Ep�/R���"2�س�sJ�U�h������������K������W���j?�M)���t�RM"F:@¤w3
��pc��$���ϑ�5�I��A:`򄠋
KHXR}�;�(ºX�ю�p���
���wC��l��@����D�Ǥ��C���Mvs`�^����{E��w�������YD��=� T�Bt�R�����x���i�J��m'�M� ���8z[�E�C���Q'��_���$F�9�h3&E̦���՚j[d��OdW���'��c� >�˭�6�R$o|��at8��wm�~IpC�i�-Y>�������4H����\�-�$�o�y����H�٤)�T�Y��������mI�N�i����Q�I}�-�х�J*�C�Ed��#+u>xgA�9��%�@R9�g��_�:b�}Eld�X�����o~X��Jfl�W���?q5aj�7�K#�� XO��\�s����S�I!��OA�$l�``�d�5.dP�������]�F�Y��!�,���bH�?wk&ؤw�q9��V�Y*"E�c��t�J�l�'6�`���vI���L�<�,s�|��Ç�Ԍ@}�1�J�UL<4tk-����C�-�+lWE�?{��'�5�R�^y��_4���/���
�T���O� �o����S'�+��R�Ϳd��/v8'`S��j�����b(=�:8���pXom�N��
7������=�1�٭�R�cԮ��Ɗ�eSe̳�y-�z��b�7�[7Ғ~�T]��T�T���F!(@����`�J���	ZAh�6k!i'�ᜈ��C�59(����J��~�&�dH�X�m�`���\�|�W�laxb4�0��2�a��5Pe`,�=ĨͶ¢�f�����؉b�k������v���0��>J>��
+� 	�q�B���ٕ�f7�:Z�G+�Z���<�.�lz�8.)��t���>C �Q؏�y:��� r���Dt~B��ւ6ȕS�Ꮬ�y���v2-�yA����O)wDmF<�rIy� x���Q��#:(�BX�|�=�iܤX���p�����t-8��Ssf����L��8F;Y0O��1�I&�/3��dx�\��Κ�t��9L$��(5 �
!��\���J�U�L;�$e����r�'��/}�o�a�W��1zZe4��n�+j�a^�(����:ߍPE���z�������%�32�#;�OK�Q��?��������A��["h��h�>�RG��q(��4D��^{�~}���7���2:0V%̡_��,��xj����~~�N �3�P	Q�Qj�a�2�]߀(+���AF���D�d&�_{��hT(�`}�W�D_ �G�n�S�Zy�����1�u��?�kt��.H�{��'��V)��%^�ࡵ�����+AZ%�%t��q����ɭ_a��G�V��QF�	�!wm�(]��׈�R��?֚��߰��s�Q!j��cĖJW�@%�sGH)��h�ۍo�؞�#N�8��DH����o��C>$I��	[�V��������H��T��l�OnN��I��惎X���3���pT���^��ޙ�(i5{���f��r���sT��mo4�|lW�����{Y<!�2>sE�7���;�x9��/~qd���Q��F6�2��t"��1�|���W����>/�=���S�-�YM3��B��#.�mM��X���벒#*��';��,�{;y"���(����o�U���@A��ԀN��.q:�����|1�j<�λ��b:�V��2#���{��G�`���)�{r{�W�|��5�Ym'��b�</�5��,%a��}�z$=80/���#;�7u���x��q.��y�K���Ӥ��1�X1V(z�MWӎr��A�`\[���	S����,�������H/`�h�盳��=��rI�EN�!��L�j��]~:(��n�J�����~��=�����y�&JA8C�t�
�?�6G�n�UǕ2"O�[��A��9�b	��7���+�[ή��-��P��k� `�3�8��=֠�TS Ap^\�j�$�U=2�����-��+NFY5,�2x��|�k�.� ��MRIɜ�1O��O�R7px��ұ��mG����)��O�ʍ��=�n����D�d�L�V����$�<UK��N.�����D��dL�-�{A~����y�X��T8�J�.O������11�������2�ң����hG��;��@+i^f�i���M��9�o3��6�J��U��es=:�N0;T)�6��� �9��ě��8dJ��m~����F��=��{���Y(<�C~���(�����Е��"c��RѥLF��71_p�^\.�'�G��l5w��d�-I�������6Y��/�Aff�!RH���tB~�P��ե��wbU�Γ�3��j
��ےiJ⫳�v���d�+"�Y����:�;;6����*��:-1�Ukd��g/|�،K[�À������m���](�+5ɉ�@rk]l�t���>�{d��d���`4!����}{~�ŖB�Ao�C�؞Ŭ%ڮVN�t��o����qt�.8��Pl&Ms�����R�5>���v��\�sňS6s��!���_ϩ�Uө�PtT-�	m�$�.+��Y| ��W�����#m������n�{�-���
�{h��ˋXmK�dì�aP�c�&��^��U�YW��"[n�>.�����>�*��l��ك<��z�yM�f
�^��7�5�Ih���^��R�X>i�T��~N����o���Ql�&.�%sS�f �|,r��x��b%��(��ܙ$��G�%�
��tB�=?�7��OC���o���yB@�>6D�m"�/�QI�+a�r0�Ijlp�R�R�\���4U �sYF#	ӏ����bC}T]��m�P(1�V �.��@r�~��ط�h+��}��)k�)x�.���	H78򼶩'��S�n�#�h}��Y��+lP?J�h��<:s���ɧ+7g~yLP��T��	m���&U�7^"�:��R�T ���1gc����w��/��E��ـ@)i6��d\�k��]JQ&�e�<O{����@ �&�
�N�Y�JM�5�݌���n����6�w��wnջr�~���o�W{G�:˃���g%�14�U�b�cq�Fo��yE�����C'��R��RK� W�s�'r	ӂ	�#~��'��Zx���3���v8#��[���]u���JL��<��z*�c��l42Ѱ���	�ٮ���4
U�{�ߦ����c�¢?�F�
���`��z�p��I/��,���;�0�h���Y̡T&"�)K͇�g/�.8H�}HDk㴲1�r9�e]�_�s�#,��=���NSuiīZ�����J�� �Ig��5�څTT���*m��Q8��A̖?�q���(�[�\�r�i�C�օH硙j$��dO:���%�c�-���t�d�&��g�lv�_�aQ�8"����^*��&7�wL�Yt|s��Rp�,��<, �.�a:HV�~Q�+��)�<o����5:�SΪ8	{G�(�����,�Ra������S�~��X�93��NCk� ���X�E8{16�
��ƞ #}]��a5M�=>���}�4"+z��"\L���Wr��mic<��� �N�ovnA��"�r�C��+L��t"M[��]���K׎"��9���R{�I3�v/���FZ�=��s��-�F!;���F��6�_&j����a�:ݭ� �j��I�n$;O,_�ba]F�H�ya�k���]����+���sb�4�6�:f�Ui����5�K�vm�qt3�Zn��_�%�$�	+Q� �ل �.,T���۰J@7��ѵ��(r�FX]Z�q�w|��\t��RW�]�z�c
��>��+�"5��e�3v�Ty�{P�֌�'	�����	m����`�e�|����e�q(�n�;3���3��0N�6X5M�I,<���>�?��V�s��Þ��Kf؀�#��ϒ�r�Gs�j<"�-�W;����������!GʫtHBh���>��!��
O�g�I��;�܊"��J:�#`6�����fU����￦�ƗL��WEZ�^��7<��!��	����x�z���f��R��)=�Ӥ�k��U�n��Bi~t��DԻ�=���!x��&�u9$�4��A0��6͏#�,$��ui�%J������0p�
�p�ڠFZ���;��F���c*��K���h:�*鎾�)j.�q�b�ޭ@🍄����G�J���S�9H�st�gЙ����,Lj��C��O��U-"AI��z�� e�o�L@��(��|v�ϼ����7=BGҩ~���o����m���K�÷�߱����Z�KY�R�TR�s,{�I���f��h�?�cj����d�3@�����i��)���+�)�_[ �8�˄��ܗ�G�ƻl��X��"�"�;k4yW��a ȍ���{� #
EF��{�(�`$l�}�?9y�^���S�jG_x.���+��k�{�	u6���zj�P�<�l�|T#W:�yU_vdW�p��KA2�V�H���4�V�r����O-��p�����z\�/��7�.����;i~���T�.�䖟#�:j<)���ۯ�V�K�?B���3�R?2@��T��J,]DeF��A���}7y�%�aRK ���O���5�"S���dZ�('�^8E�/���ȝ��aV��N�h�G�M�<�9��r\G��N/Zx	���@���g��_�=b�l	��/*�L!�5�^��	�8�=_<Zi*^�h,����έ x�:"ϩٛ��j��`F[�ly�g&�<� 1��FI1�^��X� ��2�ĳ�u8���`�h��3���IS[,K���-�����	Do|��K���ɔ�m�^�M�'�P�*���߽�o��P:	�6�ȣ9��_��a�J�T
���3q�+�NU�d��Z� ��*h2hd �B-��+}L=� ���mϷ&�r�FFX?<�j���4)�oIF�vbh�{+w��h��	
<}�l��s���n|�B�96] ��}��,[� ���&�k3 ,�n��K��C���U����d.;�Y	`��C��h�Kh�Ն���ji���A�W���zڛ	3l""!� ��xJ����e�Pէ[2ڌ%LK���
h�i,>�6*1�a��{�i��ғ�k�,��-�F �:
|�L]�ɸ��؟)�/�x	�`���#(�[s��蠯M��8ƶJ�&�~P�@���g��ڐؐ{c��R~��I�46nGs��55�1�>�=��w��g-�(j�#��	*���*�DZu���B�� �ޭV�nޗ<����u�\2��<�'n��Y��+�ь���"��G6���B��=�w��̼1���vo��%*D�4����f��"M�0	Q�0��YͰ���-{��i�T�V����}��$�(@p�t�ѡ�%]sG��W��m��M�L`��Sc�9r��m4T	h`�<3����zqz�UH�U�{Z4ȀŲN�5��vL}����M��P)�1�(k,�본:H-�}�>����J˛���`إ*˸�Y����:w&v~��U-�"5}r,��Qk�$�-�G���2�c$�B����C}~�n=�qz1T.� bJ(�ɟ�#	.âo<+ju�1���s�`�֕�t�������{�2�x���U q�~)����>U�p+�\���Jc2e4Z��\������`<xVZg4c��"��X��g�Y&PbH@@�s{�a�&�Zx���1=��;A�9Ho�:��"�e���k���b�!jy���>m��p��M�z&��JǊ���
SM����\V�[���u-�����5��S��a�#2��t7��|v����Fj�}b�p,�YkG���Ͳ����X�~|�~�8�!�Ş�>��ﻡ_������h�Or����*��uv���st��
&����@ԣCX3+B;�a��In�Dt��W��p]/fA|=+2'�j
*�u�OR��d65�Ր!��< ]%�ﴰ�*gy��O�7AS����b�[
�,�:���Ɖ����l��?���t��>���M���wYM�Kމ%݀�qP*�:h�H����d�:a��"��c"]��0�C�J��PƂp!��0��IX�j;�իJ�Ϙ2�]�Ӡ�����[tsw�6����U"d���D��w	BQ��X
^�e.a]��8x�Y�|���&G�T�����T�{��U�Z�'0��~(Rl�>,�籏/�^�6�,�Q�^Rw�2	A:O%"�%��6��W&t:$��+�o?hJ�k��x�>@Mc�D%Z5S�?�6ɺ(z��#�WF@u¡e9��z"2��4�`��yDsk��V]0�CNq�٠���U�>S��=F�������?�>�ȁJ�B�)��+��'��A�A�0&Q�x&��x1��؛�~+1Cm
|�S&���ڰUa�]�(1~p[%C���	Cv�q��W�»���(�
����W]�䨩$�����|3f`ȶ5����AD�DFòk��g!����ee�߻��8'��0i5�ݬ>P#��P�KWǉ���%Y#pw��Ҍױ(��Ba��s�i��g\���9�m�/�A�p��A9��C�19(���v��8�#Rus�F�p�B�!���lGxqس$<�O�X|_+K���-�N)�X��|HN�1��ǽ�8+������}}�4��˓;�>�2�=�3P��F4%�����d������ �EO|͠���/K 1w����y�|4�CdX��Z��!"X��ĭ]5FY+س,�f)���M m�H�*T� ����V����KǷ�r��6ԥ�R^�ꙿ*\��[gX�i�L�����^
F��n2&�c��L�}�X�b<�	�,0o�#0���!�O���̸�tJ+:m���[��'"(@�PX_+4��B$��Ki�<����sY?o�R��l�1��C��X���]u�lzȚ3�������4�6�^��]Ix��?Jk���� ��.4��x���:���չT��/<	���V|���c��A�kжXMB�Ŋ'XN�B7� �Fɑ��NUE�bZ�����O0I{*���kCb������q\-�AO��Gj��7Yl���;�#���z�WZMX?dO����?��1�g.7J6Ӝ.���c)�	��?���9����`�e3���<�y�l������'F�;��ܤy;SU�޶��!#�֤z��ox�-�܀�7m���f�[r��kT�E�j��V�Q���`.����l�	uTi�eI����,�����Џε�C֯����'�~����Q���������\�e(�̓�l�)r��x��O�R�7�~e�:��QJ�ޮ%&O�O��)�|C�4Y쌞� u�� n��*'D|�?Z�r ����0m�,�0o+ddX�*M��95^������LL{����d��҃��p��Q<ɮ�ks�����d?I�YO�\z��&|ea}�X�J�K#���y�`���Vk.O��Q������q�\��y����N�'S6I��Y�mp��Hm�8s9"yH��~�Ag`�\�8�oU�	�����o�#��s�J��(T��0}�:���i�0��B�_ֆ�>{S���|?2��h�D4E�"Rez����9�q|~�]I5���\M�Xf7R+�H��>[��@��Wi<G!���٣?�p+D.熤IY_�*'���	�xg�-� |����	��/���9g�ﰍ9"����W��_=�Eg�gy�R��_�V[��d��\9�|e.�	{���o��D�|�hz&,��Ln(z����/Δ�b⩹�%J#c�\p��vn\���?NE��^	��ri�Oc/f�R�F\ ,�FT\c���%�^m�D�c|Ɵ�/zN�o�~�K6�]偒KJ�E���+ 	���r�G�D�8��Y|�����7��g	�r~ZN�qo 0DN�ih��#Z�"�3Y)��A�Q�66�g����������4 !�P�T�h�u������c�/@�B�.���"�Ī��=�޼
yr������ )?b�mK}�`\/y�}�&���Mo����i�?�G�ƒ�)1va��I��.%�������O�<�w��jUE���d�j��h���R����η�t�ߛ�]���-4r�ܿ8�=�6��/��F�����D����}7D �N~N�q�^;z���0B����1�w�0'B)�-RM�izv�]��AQ����8W|�K�����S���z7��������tH��%�KQ_V.�A'bg�f����$��O��U�@T}|��W��"�n�)�U�[����HI���B9��{�YJ��eYl��/��".}	#>&k���⟂|�U�H>�^�lgcay�n������#��Q�y��(A�ZȯY�S��J[fٞ�i�t:ĝ�&��#��yL껐>�h�c�@gO�Y�j�A���^r�8+��I&��Q�a2�S�R���r�7\�7������}v�,���QV���Gx+W�o�;�+! *�܏��_�Z_`B�/�~'���&��P�ޛ5�m?$#+~)��5�$�*Z�L�ߎHE� 9q�^�Z��j�����f�Wv�� ޲��}H
CS�莓�.�����0f{}[�����yL�W�z�����)�O�1�{����{>�B�'�"��TI�g��]"��Q�4��oŎ�;T�NŉR���-�u�C�Y��K���P�ݔ��I�	G�*
au�����������$ř%7%���6���كf<�_'�:m��� ��>����0�SwЮ��lҪ�K��%�/��0P�ؗ;=��P�%U�l�C��%b��� �yy����Q��ޅ��c���/9%;�x�\�(�7��z�g�x!�ndN5�j�E>��3�y���2�\"�;�Vf'ah2��kSR1f{�̍�r�Sy�\�9e5�ul@X �Y��u9���|9|���Q��Fl.s!&�:��9V�>?Z��q��P�f%��~
��ۏ��%���r��`������y����%!�ћ{{8�3$٦U1=L�r���-�u�X,|e�ػ&��WA�
�*�P>������/�N�s�/����!�P�#�@t���a�&��:���scR�E���3�z��ja���[[�I�@	��+a��a@П,QbL>	���K@��+�F��S�a����=�!����,�mki2��02o~R��n����a|v�Cou�8��2c�s�Mc����^��FT"�����r���Ǝ�3!Y
O���~��lG�	ӹgφZ�2�Z�-�֮c��b{�f�;�mw�"�)s\Q�i8�"�>��騮��d���C��<^=ВuȨ��V���
�Y���9���F85|S���-�ZWc"�g�H���cyz�$Y��'��]:<la�u���Zw5�r���O�x�V�iy�?�:Z��S�A�/<O:�3t%����oi�����vʶb���\]9/� ��$�rpm��P5�= f�x��%�m*w��~Ķ���Z0��)�����	)'�(�W��D�s�_+��U���oJ=�Ϫ���0"(�U�P^� ��rz(�]((��t���㎝"$Sz��H�]ݦ&w �2AL(N�~8"ܨ�Re=<oi^�2�ӎ$͓����\��-�^$����n
��aa,[�xX��֊!Ss����n@�۲�G����Y��t�p�w���
��.���*�����m͊�H�h�P�3�f��Rs�e��՗����f�ly�H�|����mN��n�)��6���]w_�;q��'	���G7N�A�B�T��{��{[ax���g~Pl{RIZ�J5���%��f���U�����g^���W��ly�L�N��3 KIq�|��4@ 7J�u��vU���FԮ�Z���)pn�1.�Eh����Ρ�8INlR��E���6��3�0��"�MIz�z�(��VN�U��]���ǩ�E���o6���>�5���pj��Um�ߝ��
Rk��鎃x�V�zz�����Qt>�²c��X�Ԭ�B���`R����J+�
�O��kd��%*0FrE��)��t��tXxP�7:oY��\@kb�rs�Zu��h-N2�R E��Hn�d��T����ӏ�i��n[����M��/c�۝F�)R�U�A4Ҡ��vOz^@-��F���.ǝ�̂�pQ����!n�������/z0	����)��:_�,k�Cđ%��S�G�~F�?:\4���v)�ƐS��	������s �"�ر�i��=�Ǔ��ӄ�G__�]�Q��hkS��A�l�±S�LY#Y��_,-TM���X�H����R�A��Qm��g��/���8"� ꤈��C|"�TCF#��_�@ ǚ랡j�<���������>�	!���^>3'�^�d�Ə���c���o�����J?���q�Q 5�r{V~
F�u#; �ȏu�X{���_͞UGTN�O���Ԍ����õV/�z3��j�e��&Ԓ�.'��E�*�I�b���]�k�+e9��ێҐ���0�bbj5��x+4m�4�w�]�����5��+���\����9bI>^b
��	Ƣ��R�A�v	��&�*�l���v0�(�@g�7��F/�D3���q�b-�V{�
z����>���� r�E�����Q~Xc"F�^+$쳾ʭ�{�r�/f�̀��0	7�?Z��L���ӡ��A¶}Kǉ;����ҿݍ=a	��O;Fn����m�Bx�+�Ί�<����;��v�w�]|������ ��sM����T�*L|SwxsK�a�#����D�Rw�fp��Cs����F�E�ʣ_;7r�O$��@��#�K�lo�5Rˁ��U:�����Έ�6���}���x�Y�J-c�u;���C{�����v`2�n��5r�ޖ�?�Q/�?
u=�d��B'��q�C��1�����[��"Cp�/l8�/b�W+
��u�A��G�R���űɟ����KV¬UX�x�����蘔.@� �ς?�h-f��m�&�)������,�a��m��������FIޑ�T����?��X�������
�� ���=Ӣ��&9����pc�|YA�{�U���7(N�A�hy&^w���;��<��9�ʎ�x�/K��I�'�b�.x,3�K�bDg��C^s4AB�v�3�h�_�q����\�X>���Z�i&�'�9��`�	�I܎������-��+Me��告��6`�*��J{���^���h�Oc�:[�r9���Z�q|�B���jxυ�
\�e����ޏ�p;��`ޥ�3�sF��geWń�hs� 9i����9U*�[WLC�^��d�Z����[[�"��i�i
�1�b��C�3��n��l!��&�q]d�c|Pj��|B=�������(����)�����u�v�#����I����Ok�*lǋ���S��EX�]��S�� �B�7�b� ~IR�RlU���'4�dEF�����4@��%dZ�6��#��J3r�>�[S�~n�FA8����������l����	�ŭ~��1���>ĩ��m�e3�h���w����B��f�*<h��<�����#� ��q��Yr"
�&xn��T�9��x~��5�WKͅwHmNs{B�Un�g^����)�6���2Z�0�
�:��|Q�3T�;h�:�;��X���z��*B�N��UP,�NkQs�]qRF�\��╿>�:�?�`Ge��Lҡ|���?�-'�Xֱ蒕�~(��C�Km����h��J!�z�γz�O���eͪ֊���$�MZ�:�QSO:	G��'�X�]�۳Žt�2I� �%�ת�_�U�����<��AA8��Uhy��I�a���[H�L����ۢ����-K씭��Yf�4	*.]��؅�4��?T�I�҇C9�wl:t.HWw|���YC>�<MϬRaƭ���8xez<k}# ���W٦��t�D�����rs8�X��i$:����/S=$�V;�"��6���L��09D���V5j�8����{�A(7慞����G�P���F�����P��0�az�V�J�����޺�$��
k��Xۧ�B�<�\.jW����4����{t���Ll�v.|�e,�_������9S�b��ny�w��!>�N��e��%�����-��9(8�������{�S��<ѱ�AfO��'*6g�8�8́�Qf�z�:3����H�<�~��j��f_�"4ׅ�ȥ��ߒ)O�E"����Y�Z��|�z�UhY�(����3��H�S�ml�|�S�Um���0!������y��i~�Ǔd��XK��5�
��xΌ�+s�E'[��l�w3J����4���5�h�E]y}_��J��+A;G%r����0����0Y�M4h(�rGP�s��T�����}N�%�p��(+�a�ƌ}��D��|��P��tA�-������1[n�e������'�]�.\�N)�7���ħx�~�����|�����S�˫RK�X�}-}�~�� z}Y���ZG�I���^{)��<Tȝ�����1�[��M �[���l��4M<b��#����v��Q�4���U�н�3�bT����������2��(�|�s���R#<{��x�%z7v������I��<��'�x��m!!WĮ[4|�ڼ�b���O�pkװ�γ����l��:�)ݥU�'�m��/��V����/�wa�%��7-�ށP��L�S1�䓨z0���	I'M��#-��bR�'���h.#��� �;绛���4�	Ͳ��ƣ{a�3�m�jn�Vbc���7��k���PG��,#n4��5���bai%Р�WT�(���Z����n��a�^y��Pb&!�[���Ë����VCL![��K'�^��Y�x���׳�M��_m����� ;�A2���  ��n��&�0�?�`���Y��JT�%@�S`��4���}GS��툧��Y.Ѵ�r�8�]8!_�|-M_��AVm��8v���Je�/ub�Њ� ʅ9>�)���� ��:�� �p |w��a�L8�N�2�yq�X*b�U֡���P���H�ܦ�0��tKE�h~Gv��w���w��
�D�'S����\ݭ�/"�������;b�N�zY�����û���#��%}!�Yx�C�߆�(��7h͡�O�x��Q�e8��wl�)nA�7�z��"9q������ �!��[b+T��ރw��m �<�=J�1�!�u���(��Q������4���N���f	{ b��gS�r���:�hD<,�Rk�)3J�0�޲?V�9���	i�i�e������4��A� ��%1��y�_���8�Q*�$�޸�U_�%�p��X�#J����؋���)��%C��9{[�|��#�>q<�W3lB+;�WĔ/��=2�q(ɩฉLh"�u� �����g/���,�6V=t����̡Q��Ĕ\4�@�6k��L�q�g�P�%�� ��(����w�K.��*��ay'{AVj�R,U
^�1)�}�P�)lw�@�}�!�ZnYŚ`ؚߨ�X���1� �P�`��	_%�HZ��o�ː�(*�"�=.e� >n�����a�N+��T�j���2S�����������2�D�6�%���5}�&����1G�6�t�O�E��B{�Z�k�~Mwj9𼉷�:��R��}/��4rx���@��J��i�K���ɗ�M炙��X*)���������/zĺ��1?�f�:�`5�\2�!:#5|G����|3�l{���&	�J��� �9�M���9�̀Ig��Í�Od���37&o�}Xe���b���{t��n���^�a�`���(Ě�;����^q���K#�*�ޑ�W�E��)��_t`m��F��~�W�s���ӈ���j�A�;Jd�#�RR�.N�RۙD�����X�k�"#��;�I�B �h}���;~�[�6а��������B���)�p�;�{L�	h���`|�!�qp:~K�q,��	��J9!V"�X%��V*G����<� s��X?N�Q��H#�|�qc5��#�4H�'�-t��ԧm^b�i\��=�_���GGα��9q�~hg�;6�&������E�o��xs#Hx���'<aЬ�C���K9��'��Z�'���ȹ~����T�������aD�*'dqZ+͝��Nt9\���N��l�p����An��=��W�0�_�LԲϣ^9Ew�o_�|���`Nx�\65t�$VVNj��X/LvL��%�K���Z�+�GY �3�M�.a�)U�o4ɜJ��en��8Q���Ì�����g`H=����Մ��v�(9їC�Z���c�uS�mz�|�W3ލ)�q�h�FWL�^�ha��Q�ܛ�݀�y7��5�P��nK�?����؟��ۨ£��{lfM��Q�����vԱ��k'�5�p�uWG-��]�;;� p�_�}L�����b�$WH�V?!�Y�H?}�HM�@ɍ������ߡ�7R�|4�T`צ�/�	eć��,x����Ф�� oΔ�xN�&�gq���/���"��Z����Y�� ��N�g�zژ��%W��Y�|�|��	B�E@���`|�sOU�=������O �׷+U��8v�[f�]3��pe���8�ӗ�:�(J�"�Z�\8^�@?��#e�fܑ���2t�� ��3,N�{�Zs_ ��d�3�2iN�gB?3j�9�>��D���ZW��]���j�(.&:l~r����R
T3�!�J6�E�S��šfj��Qy}�����w��i�2�ʐd�ῧA�Ic;f{��_ڿ�q2��������<
G�	��/��~\��?�S��7$����D���Q�TƺӴUB"S����c���ڗ�}�,�2�18=o91����Dq6�aӵ.���s�!_Ob�Θ���u�������O����ߖ����\b��������Dy9M��.��N�+:�CT<Ĉ�J=�����Q(��D>UM�__�k+�pj��ҪVl�Lٿ�Υ����77�:�+��u��m�TD(��өu��V�]ˀ*}CK��e��R;�@Z{�Lg#Q	���`#�#�_�O�QFh�{�������p&y��ߚG`e���E?��(�v�<����'�^����2ގrD��P�F��=�?��s�rJ���{�oJr��]9��U�C!��l���I}k�RQ�3ɞ�	 _憕�B���|���xe�҆`���F��X��߷�VSu��5�0Q����[W��hhZi5b��e��(~���z8��=�/�E�8��SU�vv9�~b�L�^��f�#<e t��9-,� �]���4�Z�����B`�����.��'�a���x�`�aǓ�z��R�8_���z�2r�cW9�ꩮ�1u�+���PA�����~��l�1W��~<�����׽�س'�;�@_ml�h�;�]�|���XD���\�����]�k��CP�(�n?�kn�������p���I�4��:�Do�a���ZӚ�}�hی�\��{h��N����������P�&�{�o"lגn�����Wmm�v���I��5L�iF����l-��d,z�q�����zϢӉ�����HN�͕z�w�B�d��.��P�M��2���N�e�a��?�)�[���U��9�FdCj*��S"4!�eTs%������ְ]'�KBZ����A%#S���j�Y�E�ӛ��'��!�N�/�d���7�#MW2����GH�L25���4���I3i:`8�`��X�m,��ȿ��Ô��b;���[�Ku��]|��a��%���0�17�,o�ɏ��v\��t�]( ��;�j�ao'�S*�ak)c2�va�_�;r �
�ӯv3ˡ���mR�$�O�+ݓ���u��yLhl�1���O�-�A2�H������I�O50t�4�^nw�EQr�f�Hb{58ڍxf�>a����C�EmB�9���9Xby��Ca�,	Q+��~��<W����j��1�V�Z���������+�4�e���}�����=�|����t�" �Dlq��Ɲ�U*��M��`������N��)H��$>P8�&�z���Pt�Ux;yQ�`�~Wy����9��r!w�%8k�ޢg�*��#;�2�]�����N�?7bm�w�ON�sG��`��O�1��J�
�Ӏ�!)|�.P�]_�:a%�8�a�08 �pL�o�\~�-�C���WHGb'�qT��A��`�D�[~�BtXRɳW�c� �M�]b�� |�{9���x�C��_z ���-co�y<g�� o:��$Q�\�����Hл-��"!o����J'�E�Of	�%X{֢��7yn���Ǟ)�����,0f*��=S k�ʙ�^|���r�Gσ��O���0c�Ha}�� �r���t�
j�L��3N�DiP�(6BQ3�6L�?��E��`I�qS�/����
�fz�Y�����w���F��`�7?xi_얺>�[�������B���mc&IQx|(���L�}��G�S'���Ffa��2��Å�$�*/4�������XYoQ Of����G�?�rnJ�f�ybiQ<!9Ӫ�\�'#hɩpʴ���GZ��ɰUf��J۝GX��~$h�<��c�X���U[���[��Mv�]�v����]�g��w�֥�R7��/B�k}c!�@i�?Y	,r�B{Qf2kj<	6�	��v�$0j�
��M��/���nP�gj�!��x�.�7��VQiY�0�U�������8��Cy�b�!fX8m!�0ԝ�G�j?��[�f�E�
��,�h^�M�/�"|��Ta̱�U���댯��I�#
tچK ���4����L�g �)w��H�a�yP�ח��?��Ya��Y*4*��o����:u��3�������d��b�ϏP��M���5��&���ВD��T
/���������!�g�/?"^z��k��5(-2"��t���j������}��P�G��	]��GV���.K�!�� ������A
!���s��V�H�ǰ�<+~<��~bT�4+��r/�ـ&%�b-�k,�5!]��
�:v��k%�i��eGx������O2���5ъ��93��58�#�OI� �I`��4��x��"l���a��f:�J��Lן]�	�|df�c��u�Q¿b�|�[�(��7<���Qϣ��װ&�)�-����>/�.���c��ړhx�z)K/�:X�(�Ϗ�nt
`�K\fe2r>��<���i�Y91W�Ҡ�Rs^HC&mv�����I�3
�d��\e��`Y��i/g�e���[��]�Ҟ��T1���Z8�M���\�
���4�kt�(����^�{�d�=<i�[�����qL�i�v2u��[s-�J����_@4V=(t~��fY1Rjrb��Zu�޺��#]��ǩ���0��)�������R��4�R���5`�7S��_6$��*�L����\ކY�W��v�^��U��:����5�������L"As`Tm��<k�_�+�岞�i�Γ�C�/��OP�����4��M��	OXq��Ee���1�:�Y+��E0�qk�2�x\j���?�u2c�22��mE����#�4l:<��.��V�zS��T�bH@�l�#t�k������U� crK���G�9}�i��ˣB�;���>���U7��'k��P\��'�_��f��@���}�&X�Pc��Գ�dpg8
S������_�ӈP�C'3w���5�.��}�Bb�e�F�� ��s�S�,���n	, -can�k�������l��LX*� ĉ6��mж.(��,�ƒꕮ5��H���ܔ����Ѵ����SF�U�����%�^vґ�7>I{r&{������ur����ʟ��7���.�rDxwND��Y��-�38�Z�eM����U@*��=� �-�ч��	�}�,ɵ�B�qI�^{u����Z��T���a��.־���i�6×���x�����J�+�V��4�����8q��n�)��,P�ʒ����6��\�`�LX|����Wj�^�s�2+|�����U���q��+G_M�}!��NbP��p�M���jEb��x�� �0\t�j�RdO�����	b��]��o���8˜I1�nxw�)�o)	��ƚ�� LO�9>���_��$q�����*3���ǡ�l��y+qIK��5@�=J�rQHf*�ͅ-3q���5g9���k�_��9Ϝ�� �ƍ��b�ؑ+Vov��G�7�@P��#�݇TYY7�[�~�T��l���q�j@v껔�n��Ϯ��uva�H)����7t}���^��_(���q���*m��S��r�rk=0ہ�s¸��Y�ݡ'��`Ӻ�!z�/')ꎒ�o��e�Bv%���CcF��1���XJa��?x5ڇ��cx��v�63E�DZ:y�����d����.wx%?�>'7�t#,l,`@�����l�<�#�yC��_2ם�frWg�������^����^���@=W'Vvm� LA���뇳+h�Q�_��)'�Ǘ�5:�!��c�Ϫx��/��,F�.�5	�j!�c7���s��)�}D,�(x���N�k{'�{BeS㼟��.1D
��\�&�[Ѡ�����.j"G��^�F1C�Ʒ��+9�6���v����(F?��ʬ�K{��zĂ삧��g�$J漙G���곊f���	�#���q�:�Ɓ�/�A����BV�/��������g�G.�����9+g�t��cdQ��)�����T>ؾ��h[�i>�����-B�;��fg�#��_K���3�k�_[�uϺrS
"�[���4J�=�'�l*�w�}�(�i8��ɜ>[{���$7�9�m�mt�5�Z^��e}��u�4��0����Ҵw��UnT,� .��*)�yK�賿Z���w�4d��k!�Lf3�`��U���B�1<�W ��O��#��8��;s~M�M�q�������}A�k(�~���dt���W�T.�Y<�*���>x��Uk8�`\8��זe0����l0��(m*Q֖.Ǒ��w[<�x����_?�3Y�������¤��~���Κ����� G9�Z��P<��w,>�pJ�8�2�n��4vFF�W1�zT�tje�k��H{�i��PQ��A�hSBĊv�]��կ��*y�.m`�e}�#+k���c�����IVPM*��.GUW_W$m>�=���u�g�v� ����)V��
h���n��N⑅P��.�� *=�mZ�y�3|��w"\�8��&���(Ч�`C�Y��Y9ٟ(�h��@�މ���Y4���<�������Qy:�EiN8-����(Z��i���~�Ƶ��q�4h[��~�D'f]���95�!�.�;��~��
u+�n/��
��R~b��ՙ1^�}�T�Bl�=Cl�O�[�l\IS�=�&�빁��n���ȇ���6k7���b���3��)��+�<Y�tM-i	��^�nU�Ie�F�l@e��񾏺(�p_�)��ɶ|N[�a���N�N"Gx��#)9����Df4�`�&O>^'��r�!u�fZ&����`���r�rp5�S&���W�՝�茏	x�mk|ܽƤ/�T}�5��bl�3�4��0����VG��|GQ�Nc����SjnO�\���AJ����n���N��g^�������@\r����6 �ņf��d�A�S��W�(8�o�ǥqIf	}��@_=5�z=�T����1,c��;���۶����Ӥ�q��`N'_�Kz/A�\��N+5�߉��kC4�:��0m��h�Н�b�:���6`�8�Ei�y�J�/o#T�oP�V��Dp�h�f��2QU��jj������=�f���g*_HXu-�}��$M꩙g�Jd�+`�Duo�ƀ���2����-1�W6�@ƪ�xN��R�J��&k��(�ժWڂs�'O���_��7�o���s�"���n���Y�_����U%.���M�n7�Hc�
Jv�%�ҝ���#�1�膝 �vA�� @�"�a�^-��U<Y�%,X|r$U �:�`K3����p�T�_a����F����O�u����4Ns 	�~HN���J�i�ʰ�v/׭��t�՜�n�ȎJW��tTf�UB�%�X� )�Tج�E9|(�X|�@:���G��X�^y��ʛd��8Ms�z9<E�B�cQ��roҤa"ɔT&��m�<�vJ�^���)���Y�;�B�Ra��̈́}2B�f��L ��ɏ���~�eL������9Ȝ_iwrZ&F���az� r-�]S�����j�`X�|�1=r��r���G|j���k���K4}rZ�D_&����ձ�	t��B�� _��܌��J�1"O���"���R�p��(��-T5� _��61�ڎ�?����3��A�aX�x�N�==���-��;�W�J	o��g�q��D����Qף���Q6�w,4 F��@��H6LP*�J�"�-��R ��ſ�x������=���$�nvt�.!�)Q?6!�M>c�"s�)y�x����P�����|������U�О�>DRX$�P`^�<��з��S��l,PR�p'b2>��Ai�[��p���K�|����(�T����`��6
�P7 -���xg��)N��.�y����g͐>�^ЛY�e�^�&�Bc˭��$��2A�Eb���`2W�IP��z�}�6x��F��2����������3�u�C��i�-��aIsX���	Q=Gq]�$J(�p�P�� `_��n/J$aGNY�F͖_�8$t�M�EF0�T\��19�wC�����0��f�(&<o��i�|���˵�i i�JF�����{8n��o���L��*��p���"�G��t�N���$���b�	�>քT���,q+jEh2]6B�7�qLޜ9M�eQ���틡~Dϙ����|�R�"�I�{ �َ%��ZO�j͖;�=�끊yl�V��p�{�,�G��^˯�- ��"��ZCџwx�W��t�ԓ�915i�S��f�;���X�d�=w&_�U7xKT�g�c2�vy��"�D�k�a|3�_KJX�"����dsG���p���f�6��#�o��}�s�RNGM\���PY�A⟻X!ߋW�DڥQ��lq}�K�w�Qک���uɞ8�f�7H��bH�SY���I	�G�p,���w��eI�O�S��v,T+�/��M���%_*(�1S������G�!k�
T�J�U�z�l|�oKt�L�ޫU��7We���C ������:�W�^%r�~$]m�Z��4����+�����T�K	�]���9��&	:qcFh�O���,�_ekl��Zb���Yqa��X�m�B�*;���z�{�~���rn?L���I^3��u9�tg}���^�k'
����=�̓�fV
�.�	p��a_ᄛl'<�I��a/�3�bԈ�t��]~G@=ұv!\�t�b��M�e�- �5�&�ԳV"�]����>c�ki��A���A:`�UE�=l&C�+`B��8�b�x�5�܋��P���፼�yT���"����垨ـ1
{*����[v�N�
j����]G��ώ1J�� ��?P42u=�9kVg7�RM6�^���S5���z

�&�g��O�4�c��x���7(�oV��a���U:W��2.D�W��v�����e������GHM0�g9;[pm�PhHB�����V����hkd*��ܮ�%A�"�BW�)l�u�6�0s9;�p�5Y�u�y�\U��x��zS���I��)�r7��%-l�m��&4����9f߮�ȼ����b!ΩA�}w��?i�ɑ�6c�N�W3۳�ۤq���ƹ���ްʐٔ�A�z�0�%FH�N)ܧpF��|F�0+���#�e�| �D�H�ب�����ł��W>`=Il�׻�����t,4w�)�m\_�������;��%Xk3�ʵ�r �ɺ���J����x`+�#l�םvj�E(�,iA%����.=q���Y1�rk@�o����E��LZ�v�nL�S�_?�㤃Ӌ��b�(@;Ss���y�`�|C�l<?ב��>Yړ�0ە�o�] ϣ�6�i/���T0A��Š/���)�&�y%��J��qb �X�x�'G1��a �x���)�f����޻H
k�R�r���x��3���TH�!��7A@��0����}0�;��'�-�j��Q�ᷬ�z�opp�8�YIqG3X�VT�%�)��D��#��,�Q�����
x����L��c��zq��;��� �i`��Kɓ��߲��]c�A��2A��W�FD]��ɞ��҄�u� �O��t�
�gX��a`������KC�=E���c�9-�)��%���$��F\ji��i�Y�7��v6;�4AF�p����_�P����b��V��6R�����ѝ���1hWL\�^u� �N�
��a�$me�Ԓ�����K�uw�
�I����:H0&j��o+DP&�8��~�DofJ��@=�Y��]W�L��KJ׹6L;>x[d�Yg���ı~��ŖKe�h��X���K��C�zh��^<��L�2E�ӄ]�������c��Ͼ�w�tR����4?Jo���,~��9�t�7�5�]�� �C�Q"PD�=_�ˊ(�A�]�z�+�5��2�G�B��٦ ?��G�������^���� �L e.�B�}3U60u8g)���,�/��U[�nm}79D}xq�kM��R�u�ڎ���j�C�}�������|�G7��؍�!���}�F�6���7����̇Sq��b\y=��$�B�z��\/P׺��/�Xvޒ�{(�WU�ψ���`���Nº�{v�s�����{�ڨ6Lu��v�J�a@ҘP��2�v�����j����=�l��(��%���,��]�_�ʑ�ǱJI��W�D���Օ�fZd�s�mv�%I�P�Kj���\)���I�>�g���䝽�A���Z�\��#CƐ��Q� ��x2����y̚h'�$���q&#Xq؝�W(W&r�p�0K�"��H��?��/ja�,�W7�*A/��Ӑ?@��63��8��SQKY�il�����z�|K��M M_7 ��%�m&M�˚�9FS1� �"�$l�G��_���MM��V��?!��q�[Y�c�b���tzF���9[m��O�K��J�U���F��yC�Hl��m�g�X���~�	���f�aQ}�b�+<
��,�IШ�5F����
� ��)�8=�L�:�J|Y{6B-�4���ȇ�_2��ת�����O;͏�n���I8o�5M����v��T?"���!ԩ���~�B�oE�M�[�= �>�L��i��6�L�A覕�N5��?��ݻ ��е$a"���o�7�G:ڦ�ekFl�;,Bh&�[��}��s�O!:u�
�SdP�E�/k**䞢����8k���,M��df�U/
���xF�w38���ϻ�l�M�A���㊛�^��+n*`��4g#�_�M���؇̆���9�;-�Xk�LыG������V���X^ngv~l=���x/h�q�k<C����9�a��;�*u����^f�Ņ�5~�l?ϺVfuxq�W��I���×�3Ԉ��,mr�/ :�o�����"P+���g>)ҫ�Y��Y�p?��h��1����i
��N�H� �J	���@mۏ��
u������ah��!��Qa��`�XGm�/���7��JQYz?�����Å%[�
�x+�)@2/�8�sN�L5��S�^��ٯ{�R0դ����Cgvm'�h�|<V4 �t�iʀ=H&�d9��y�'���XwD�{��Gds�擼����ӓ��}��3v�+�'��K��H��˨�Ak����C���~�?9���!�7շp�Ub�O[֮�3��Jb�đ��:���|�3`�J!Ԗ�`m@z�zA�L��ӊʘiBh�6�Q�*?��K�ψ�q���Ǘ���1d}���0��t��m�i�CL�u�Cu1��%Ì�`ݚx-D�.T��σ��alnv�*�DۍHB�ՙl�07z�m"�ʚ�Y�����m��8ׂV/���+��I�g}S�Ω�GD[��Pс�˛Y/�`��u~�P<1{�n��&�Λh��S�Aը�.�s�i�|r���ƞ����(}�cH/�Q���y��7��?�X��V��1�d<�jg�
� <��YQ^4��U�;V�i2
������RO����C�����Y���.cT7��Ҷs��Ȳ;L�4P�F�{K�
w8� �Qp"��}�{x��N�~�l}'%MN���5�ǁ��w�=�0��)�ȷW�?�:�beXT���e�yX �$�3gxi���o�{H��1�(+THz�1����9��q�D8̉�d$4�V��^���R_�
_^:�,�Է��:����!������^�5`�8�_�VQ�C�1����.y8��i���a�9�\��"���H-�?��<�lI�_)�TU~'E%}�
�F�J4]���pz#�L=��"{a;��)D�rQd���'��������IP���9$ܢtv/Y!�ش5|w������sG��N��1{�n���ODW���o�Jy�"�[����/M���h�&u�S�;P>/l�`� ?��!�7L|��	��bg���@�a�v���\������b�#U��h�8��\$�w&@W�Hnm�S(hW-"T�z(�\�a�u��M�m`\�6��z|mb��(�qвz�>߶����ߒ�^��VS�x�3[>��� �"e6Ux'���{�U��	�U�mu���-1���Ău�T��
�W 1�x�ӟ�[�_��/�&�^���љ��.�T6�������/4���1�m*^�^��2��T)Z����(�T�֓��㉶L+8��ԛ����\�6Mw�)�SkP,+Lu�S�Q��
Ű[kdRi�m��6b���+�-$@��881ɳ����G���$U�
����T���B���2�#`St=@�%����y� G���7��Ol�r��Tk��k#�A8
gڍ�C�[��EjcUbE��V��a:�N�y�i-<X�Gd�x�������s����?�}=zz�@"!��R�'#��:����h��4��z�`���GI�A�<)9�F�32�X��Pz�k� �3�p����s��t���w#�E�I��" l|>�5�>����Q�Ϲ�0��Xu�mœ�'�&�4m�$>J���c���?s v5�Xo��&}�P�ʑ�N��G,8�_M?(�a�F ��ײ��YD��P+H��
������� �@꘺Wƭ��}T��"p`R'�1w�dF��/�(�\�[�5d(+�y�h�H�,��=\r�부���Z��5d7�8;����By�lF�au�+�r�tA�tt��C݌z��}�(�p{[2�1�^B21��s�W�sg���9�:�ӷ�Z�]��׷yc3���,���|��o�����l��o�nv�5�R��J���$ړ���F�� ����J�Q���[|y�e�@�z!�3Pr�_h'm8zn�s��ѫW�m�H i���**;��Yp�e��������5N���%�qzKL��u��u,,�e��F��FH�u�_����a�{�x7���#�zв�P.J�^c\��ք���ѯx4��3�H��a��(�5�y�YNx�Q�	�rZ��F�Ң�r9 �O�3�T������l�iS��t��{�}(R<�ݵMm�F�����5���9��=3Dʒ��c�q�9���ś�c=���P�n�	�
IȪ;\f½*"lg�i"�҅��+����܄Zq! F��R� 2�����℄A���q��#�moH�������P��	����7�!la�=[�p��\�]mnk���+��,����W��ER�����w���#*�pc��/�p�mvz2���9X�w���8�w?	&�^��Ȗ���)�����VV�b��!d�C�� �C���v��� >!�Q�TV��,ŷ�_EI�����<�l?��
_Sb����P4���{�n��$6:�HM݊�TO7���_T�ߖ���,�:9��9�Ǌ��1R�n����R��&��8/Xa�#���+���s��*GT�,U��Z<;�b��+"�����*F�Ȫ����qj�x �Zo�\�7|7�W�� �ګ��ٜ^���_5����4��M�D��hZ��B�ӮlG���Q�x`��{u$� ��\+���4�h'9ݯ�b^ۤN�n�
N���%�b�^H&��k�¬�{�2���e����4'-�s�q�g��Y�AYk������,�4��8�d3�O�Zy�������M�|��+�U�eF6HX�b��4`V?b���Ԟ�Z��\��b�����]֮����>���k)��Vܛ�;#��PxZ�w��ѕ�� �Z<��̕�"��:�zxm��I���m��=g�����8��{d-ː�G���OK���+���ðT9��@��C�&	BN�2�C	m�Ѝt�a�%)>���4���7��@��7��r�T��T�hQ�%�~���@(F��P��^2������{�&���o����ˌ��Ƿfy "�h��C!��g�U�+�����^�I#;�4O(�X�"��_�b��eY#a�-yI��)����d���
T�l��ǟ�'Y��h*��:
�n#$�e8ÿ���0KB*���+_���Q.�T`�ާ-:K��$��7�h���9h�+a�C�"$|xUs���9�~�]��J����E�����>�^����c!2���ܢ����AR~[��Ć�O%���U�Z�-`���HƏ+�4�ۓ�B���קVD�|��~,K�F���{v��|��)��+�)k�8��y=q�FRK(�c����$6��2DB'a�dϰ�ӛ=�\��J'ꔌ>c^(�S"�����ܟ�͹7���7f��>6��&s��kg����x���0���|����� A0� ��q}b"�	��ĕ��"�Gmʹ�jGJ�ϔ�B�m�!�!?����p������!�#L��/h-���ݵv+�9�!�ϼ���V�\C{��F� ,��b���������5`y��\�*�T�i��E���y,�c�*�F�����TI�2�����iS��`��#��Ԅ�K�[���n�m[�����I�BY3�����_m�V)����҂�DW�M�!k�6�.�tp�à9�8VQ
�0�'<����_攒�5�P	|�a���[ͷ"_�FS̓��``_�.�n�MY�Q�/��YW��8Hđ 9A��Y�q٪�ޥv��������A
�^��!� LkMfE����MBr��N���t�"���u��l�50Q��
x�m�1)$KxG�I7<��m9a�w�w-(1��{yj@�z�����|�z��t��^�01o60��W�!�?�;:Of�٬,JȆW�����D��u�hQ.m���ұ�AiR1.э^o���^!�N�h����
?�a�hDR�s��aи�n��)���{��(F:��=�\��n�2&�玫Eu8ʔ��1X�&��a�	�%|�u���I�yV*��՘M�$<�����{m��̓�*�7q	Y�δ�=!��Z�$�#�3K�j���\{su��RA�,x 	05��h/�G��Z�L("5DV_�Z����+��'��8�E�͠�v8��NO��"K4A����L}kk8�&��>��h�[%�����- =[:dԅ-��I��P0�P�}��?��漢��jfz�����n�xR�9���$3>Z���"��u�jlK�=�
�7���]���m����@���|B�
��y�~�����^_�*�R�r�����$��"���K�_p��v��T�mٯ�hĠ*E��(�JN���Ц�)2��ZK�*H|��)
�03���.������9>do�9�İit$R`�W��:�ݔ"/87X��~9�e�nW�v`[�Ηt@k|��8�A#�%�wF�,�5��)�j�^�M�~�zK�s%�^�}��X{/&*7ME�6�-f�#����9gv�Y��>�u���,H��Z2Û��%���@�<��ޱ��B�'	f��А��E�k��u��^�����	��vj0�9�)b���G�*�m�Z�����iO���P��	���ʫ쇳�	�Z��Q�{�p�� '�+��������2���꾖��d��"��h ��O��3$sZa?-��0������BK�+4��`��0�H��@t2b��7N*����)fu��=|��HZ��0�Rj�<���&�>^̏��>Z�;7MTVD����z��g���fe��\�D�>}�b7�FN����ʊ{֟�BX�0���$XQ.s;&�࢈ 	��ܵ���4����k;�G�c,T]��K��2�d~x�#�n��L��a��V O+�"�7p�sS���QL�_���ms�~d	}���.���붟iG����8���XbT���0�V��>,�A��H��2_�\�N2�P9�$0�r0�+h̀��[0UKB���|�kF��Eɇ�x7�]���3
�6���oN��2U��sbY���08�l!逨X�����l�.�=*z�
O�q��]���\2ϊ\Ս$� �B��� ���v�ѥ�hy�}dU���Bom蕉��9�z�3k�8�]��+�Ɲ�q�͐XRp��Z����i�Vos�}cS���z2����O�h�H��Pb�v������%>��=o�A��$=��$��:iC���� �Ώ��w��6WR�;~5ʌ���*T|Q�5��_����z�+��oy����64���=F�pESW���ho3��.t�F�hG�H8A0.ڲc6�a"�������/c�%���l1M����7��H�)���B�*K����M#_���];�I����$��q��p������l�Ҋ+ �})���d��!Yq��J��Kr���;䝠��"���q"/håN�L)�a���%�/|���w�UV4��;�6�r3�=훃��+���k�Ui}G?��Í ���ܟm2��P���`��w	��M�<�Ԥ"4�xVPg3�ޖ	��Λ�)�!)��[��I�/=כ7��ʲ�Ym��&�:��,�(:���u�J�d�V/;I]~��V3_��T��@���1�=%���G`�⭘��r)6���s÷��Ȏqx�=��zR#��A�ۢ�	:eڷ�B���c��Mkz.�VSN�������/̅�klQ뭆� d��i�O\I�3��'���ľ��� �s�Vք=��GP�@�y�_C~�M��lmys�н! i��-��8⊁X������Y�-`�=�hd_<&Y�I*��@1��Lf� mC��K��ɛ�cx�峸L��;�Y)��|;��A����7Q|��e(���^x.�\$�*����J0���R�D��'B�?ͮ��A`����a2�R���k��9ݗ��#�~߽��͛�]\ИT|/+
$`��XIH�o�ݟ�����_�����n���Ge�����⛻������w!��J��.9�$Bc�y��o��&�����Մ"�h��	�����S�i��]ݱ��B�b�	�!�NJ�������۶K��Zm4Vp�P|��-���i.���jk1�͢��1�&��N�������C���W� �2��@H��y喰53������H�J?<m�%F�pƁ��<A�Bq5-nh"zN� �+~�,���2�����bI����ۃ��"�g��a��Į��yߢ��O	�٠���A;��I�BqyB!Fd� ��U B�#F6��=�{`B��İ-i
���y*��\c�MVW��e��(Pe;���c���ƶ�z��k�Jc)�i�e=�ʿ�	=�4�d�>e�Ӊ�eqXIA�yP�N�#TD�Z��C{-�>��"l
`�#�4����#pvh�J�c���:jA���쓢�Z����E�e���M#���;��ƣ�x �NA4��l%Yb��ĳmA�����;4�t1 M����b��FO���'v7pB�m/0d)ܲ��o�mG<�����J�3H�G,̇1��O#?���t�t���F�m�������M(=�6xZL��j�n���(� C�����d=��$]�g1u��}��~E�qZe~�6a��1	�ܿ�{3��9��Ahy�+u_ZA�c��.q�6j��Ǎ�nW�=�m��s���+�l���Z�8�8�� �'�I����R2��ea�HŘ�Q6ԜŖk�׋�5 k|�p�����|��$��9^!���~c=h�T��/_����E0O鈘]-�)�Q��G���}x��S��fq"���m�ڈ��|��xC��ljw��-Y5�1�:$�v9�9����ǩӌ�����lmSeD"8��hŅ���Nk�V˰��T��AOYF�#w�V`�R.c˰�1������G��c�,���v����Z�JD���"��M7�+�;<1 �9I��F�pĎ���(Z`�������Nb}K��2	��P�v�ir�vFr7�η���>iu8?�P�%|�N�JC��*2��a�[���c{�ܩ�s���*�P�ft�#5⹈=Lَ��D`��;ª��޹�>
!O��4�y/�ͩ�
}/�x����@�$�G�Rߖ��1��ѹ�8�
�{u^v��xق�D��.?O1�lM+>��Z�����	r9�|�w��P�r�i
;��y%��c�S:�&�J�s�r5��j^`p�Oy�=�����ݖ��A��\���@ri�wI=r���'P�D�WŐ�ӑ�o��Ľ(�/F�V瑮x-���1.�,���/o/.�1V���UE�x:�#����>pQ���ķ>��)��Nf�H�i��D��S:d[_Wh��Cޔ��}��Y��6�������^���8�Y<F@ό��[㊿����L:�b���h)�Ѕ��V7R�����EH�U��E3�ֳB`��xYTT���0�5]R�{a=f6�x���B�c-�b�������|D	�����xy.��|Q��α��w�*��V��Mx	�1�e}����{�M�?���^��u~�S�s��l-^���j��-o�w�w1�!gNS.����=�<:����1ha#s��3�,GW��|^�~���b숁0/��w.���Jq���3�ڷ���;S�e�S����v
�ۮ���~g��e��A'�s�c��@0��X]���v�6�g���tQT�KX�����"-�q6�,H�Mb�c�_KXVW�L-fh0;��2wx���K�e�aNq��Gu4<��H�z6@����h�W�*�ܛLm)m����YP��Kjф�R����^���A�uJ���8%���&8i�=����7��޽C���ɝϿ��})��nST�P���]Cd�k��HD�]�(_:�k�N�����(�8
u�1�N�	X�j�e~h�����T4��G��@���+cy�2B}r�*�3_-����#����M���v�+C�Ԑ����/m��#?*�,���6O���r'�j|=Z]7�����e�.H�W��h$�[��a���HČ�׉�%�~����$&��6d�x�����f�ެU,J��1�@��7w�t.�]��{���p�?j1�@w�� \��~�1����%��y�(�J����V>��δ�;N{����?2�\(�(��G�W,���JCf����w����r&I]�̲���K�'�������k�ʈvէ�9�I��*�L��Mۋ�r�%Z7V�)�	r��4Y�7)�>�=O&s1x�t�\0����Ɯh0:�U�O�*�6
��օ��W�*���o�e�(��=˶�=���W���k{�1��#8�EA�����ELHˌ���
<��) r/�ZbۂT+N��gF��h�5�^�ѓ[�vD�/$��ݷߍ%��챆I�e����_&P�L�m^)���B��� ��	���q�E{��H����.�������d�	�䛝>L�_�T���0L�.����eI!Y���׫�P�|�!śc�JA�hE��1Y�ҷ�?��+U&=��N}lW۪��]��D�����Ę���\�9���f��i�>��|���#�-͎aT�S	���b��{ζ���vdf~Fl���lB���?dۦ�<�X=s�0ҫG:�]3e���:F����~��xT���Aa����+�u1�m�'�t2jr3ԟ?[���&o��d��h ,З���KAaW�6%þ�1 G�aP�rJ�		�׎�oE7��>��)�=�XҸe�_pG���Z��z��$$Ohn��1��|��������H�s�Һί���~<^�>�Q��A&��m����@^F&� Ԏ��Z��o9��%AD2���qtZ�K�I.2'��|&״fŌ�G��������1��>���#-��k�`
�(R��!m�7��D':��)�Y>9��
��ƹ���H�5g�1%$)=���U�Z���i�{������"�Z����k��j�t�*pIF��
Nb�����=
����]P�-�w�6�w&�[o«¨�"�����L��Ȥ��)_u��SU-�n�����ֳ8WA��F�L����Pef�������X�����~ٖиi��R�*�[z.�ΞRK������D�PA��F#3s3������h$�a��L��<�Ѧ�.�n������O��"��xA9*X�Q���yq~FTEh �2��h{uy g�8�>�B1���ru�l���q����5Za�'�$R�2�u�=��q�U�'ß=@����0��^:��#�b+���sY�J���dmLDh�Q�1m<�q��\'��������u,
��.ǽ2��ⷠ ����(�&٣�F�:�w
�C&�P{CRPg�.��cή����J��U#��{2k&z*t҆��<��*���h����~w�h1�π4=�\-���}��M~�OԉO���VB��0���*t�.
~�B��͗q���LK9"@j'�e���o��౎�JOm�n�=^U)�y��ɯv,M	�crh��&�6Kq��HCϸ�e�i�Q8�BN�*��SYd:�{)�a�'��Ӽ���b5�Z� ��m��FyPT��]J������*����r����W=&b?ViH�T�W9�����sjƅ�60�Z�)iRm�y���甏;�҈1I������D�3K�ڙ�}0���j=�Ȭ՚���Rz:�sd2�-]ʢD�Azn3�&<���"�ր0�O$=�Q���
z�r(��j���o�~�6�����da3� �'��.n���1���m7�Y�!�|H�g�Q�����$@0;���\4|Z��r!^dǸ�F��镓б0�f��-l�-�,�
h��˕����z�֨N^Mƹ>��f�"�3(���o�G�]�Qvl	W�a�57�BG	��|��
8+��|�~�}�o��i�����,�����^��RCF��ex?��7��͸��-��P�#��B�ڛ-�ۋ�f|OYp:����z��t���〩3m�b�P��qN+@%����]�>�>�=��@A⨯I!��ˎv�BѾ�Y�JE&��=r��h�v����n�/�z<y�@��sy���S���(��Pl��;��5�Z��F���1l�@��`��q��|ҕ`i㔁�Px#��T��ί����Z� �����ש�t���v�|P���Щ ^,�ӦA2E�Zd(ڬ��ẔP�Ľ�>`��!�M�6M߽e���R��/���g��E�;X~�#~)�Zٜ%ى��	:f� .�k�d��?���ԋw�z~"k����k��S�q��D7�fY����Z������J-���$U�,�l����B�!���Jd~%xB�LG��Jc����]�[4_�2�g?&��28��[�F�h�5���3yz0}(�����Y�k@ ���� �����n�fA�%���OI�c�o��������TZEOӮa��%�v�d�O�㹄R���	�lm˱3.D5Dͭ��`��"1J���#e�>>�#ߓ�(
���������YBg�\�B'���"e� ��-�~�F�l�P��:��/|P��ۥ�]}���t?�� �jn߭��ц'9��[��E�x�VK�˸Ct��T�~;�����\^G��x]����E\��E���d����bKT�%�<���&��0�>9��Yl��W��Q��?�,Џ"�����Ka���O�.�q$��IRʅfR�P��S}���됻� F�)ߐR^ޘ��W�*���N�?L�^�����Kۘe���qf	p��)*�]�o�ȭ�2q >��R�=�W������C��r�Ұ� b��_��������5���2b�Ʃ\Zy���y�O�A�u��������~�Ç�r�	j ȏ�%*Zqwb)�
���1i����3��ɮ!��Ez��Q�o��X�9/h4�s�f�5�f(�hZ�Th��a� �Nn����i�����6'k[�������H��[�-����Yzx��1u|x�p�5������=�0^����;�uϜ+[u>A��\܈��R�t���D�[i���?�D�!F�a�jv�.���^��58��N�$���z�n숑<���*�{o?<:Bۉ�&	G���cjޜ;HVBEܬƄ�`v���=��	�[�D�?�i��!��A~ͫ��VU-kY��g��.�S�2[	V#��A�L�Oj��ϯ�32�e7I��Ĵߗ����ˊ�/j:��.����2H��ը��15!�^FR�N���9�>�!�椈���e Z�I���S+0�	�;-�ַ�%�����D@Oi�j�N����*�a��F������Y<ˎ�ҽ4���=�A�����	�{�&Ib�^}����^�ZD��Y�X��ȯ�w�pښ=�V�&3)�6�6��F�ǂ��_��v��6�L%����cJeQ��2�g�>!_�P�˸�	
��*Ş���ܮ�+7�d9S�g�U�;���\st*�2M6�8�x�"W��!ڱ}#�W�8����y)"3h�8E����~,�dP0��KB�g�@mS�&�*G��|������.읝��V��̶5�N��aIFgy��̀�}��P���b�
��XK,lQ��-ek��_��U�<Ko��n8�C/ZSʘc���u>�0~��~�I߀�����ɬ��ޘ��h�jX�E}y.�ܘ�W�H�������?� ɏ3@(l���o|ðH�З�J}����̛>*o�u�pW,U?�ȕ���xw!�ӓ[���tZ3�we�g����� -�D;���h�
�-��/�}����ŗ�l�S_"��,�~���U��P��逳�򁃧r�����Y��g�u��Q�c�y���+S�%�c.��`��Ѿ[:!���_C= wO&��i���+�γ���]���vy��L�{ap�,ӳR-��M�֨e �G9��yl��� Ł�rS 6l��ǐ�D�G�����>7�����5��'���r�D�C~6���������`ռߐ�Bϔ�CvY�_�%u�) h3A���5j1@���p"ݙ$[��J��z���ŕ�:�b������V��� P���Q�J�=Gn��h�/ݑ�W��K$��X[��B
l�:1����aFo3�+�h���R܉멁y��VKl/���Ԝ�Ү�r�8?���[t�I�g�J����>{nXnz����4.�Kth�v���f�T:'�6����8���[��	���S��fGW�J"O�"S��e��B�	w˘a�Fw,��q���Bp�W�tI3D�W-����^j�MR�^W�ǰ	`��.2 � ���S�B�f.�ge�*,\��6�>��!�6N���]��G<�L�Rx#�����~Vd�'���
�ˀ�wx���q���.s��jʝre�a2|a1i��0[ݑ�c ���.���V��Y���8��q�Y�v,�\��$��
��@>��,gp�փTڏ�\�q�u�Pqݍ�E�s9gH�����#}�ޔWҨ]q��[��&��B�O�a:��c�گ��F��	A��-��Q�z!C}�����[V������"�ar"����
�-<sπ�~"/���b}��g��d�3�S�1�g��zL?��E8.�̷�w�+8�\�$G�ޥ�]�,�Nb�a}j�����G\u5B���p�uT/̺�]G�jLa@Τm�B��L���#�`�_=(T�9��(���Zj�}aս xP/L�L��\]�*,2���Q���6�E��Ǩ��I�Cd�^$~��1�U�|��+d��n���h�/�؈���}mL�_�6^�W�Q]�X;���3-�Z[�M|Ox�()i�Z��S1T��̲�~C�RY�_L /U��t/�_-��>׷)�4Ǫ��.�p�V͉.�V,�����9AO6	<�q؛v�,�{?���c�Nna �@��p��y��P��ܭ<6��Ħ��LHx���3#��"�6�a羏���а|�s�uvS��&ɱ�/oǿy��'��2�]��Ks舜��6�&�u�M
^������G.�3^8�`,g�Imd�Z�$Y��T�-�f�:��]:ThgC��|�N��A7�L�ȇ(-�Cp� 6��̐=Ʊv,�s������V�W̅�y���2�˖P�qh��7҃:Q	���w5�L�k��Ƌd�f�@V-B �|-['ݡ�8�-�ҝ'��1:K���������\��t���F��H�@���}x,yO�(��e���j;��é$���)���#_\w�f���=��M�jH.��24�F�&��'V��>\/R�x��U䨎��o�r�b�����w_&ʄ3tK[�|�2�'��pᚆ�R 5�U�u��K6Y���ɣJ�J%�E�U�q���������ֆ��3�,D �j}K��7�w���&JV���b���h�X�m5S�34J��<�e��IM-�JH�q"�f�A�gwZ�Z3�P�.�v�:ѥ�q��^PS�S΍6��b�� ��a�x!�p^��-I��=�-�~�7�����	_w�%���0!x�'�rp�zu|��w*(x�	��}n�_h@e�z�ɱ��F6s52�#�=��D$u��c�z���ɡۋ��� ����1�%��NLۚ]��@��BX���گ�h�y�����	��9D�Z�j�t��^�dv�sӼ�c�6��G��M�F��h?���oL�����U8K�͉�=7Y����D�f �EA�iM,��o��m��& ��0:���%��ϋ7�����'���{v#3���faf��v�V��f�8W�(n�ʮ�&���%��g�m��Q��`z9C�?�O�%��S�#'� .�̌s)��]s�r��0g��1�j�Y�9���Fn���I�Ԋ���G0dr d	������&����+���]3Mg�����d[������2��Lt2����=�'l|v�)�hL���W>��OT�E�'�LC����l�\f�3�����#���3���F���&Ca�
^��%jyD��V��ió�W�̺v����X������*�� D�k�IM
kTbI�U�[k�������;Wr�{#+�>j��{�-�	߳nS�6����G_��)�3�K��p�7�p\��c��.�����O����J��7���*1䥁�ɛ�B�� QV��������(1\�dH�X�r����>������]��'�2��G�Q'�o뺢�k�}�����br�f��> Q��T.H�膬l�/,��l*J������iظ��Q�Jo:��s�	ئa�W�	��'���=�(��w�f����D:7xE�E��AoI����(��j����;� O$5���֚��Ƒ��)־t?%Q��ű��
Lj�Uv�0�Ղ��@kGx�7�`hV	��H*���i��
$|!��:ݲ�[�o�FWp�_<u���#�sQ���*��	���Qrq{��v��������U�؞�!𗅆6��^�%~�V�L�������re�wC$ E34σ��k����iJ�UC�L�p��*^\��p�L��]�����yvj1�����T���Ec��j�SC�w��^��;��\��Te"� �A�'��YL�qH�V�q�F�:�_�
��Nnł���^jS1�O0n(�l�-aM܍�
2�&��q�h�$�qC�&�z�|��iŏ!q�����b_R2��g��[���9[r�X�b�ȫ OM=��%10�{�T��|_��a�ۋBO�� k�ԌN�5�8WK	���D�Q�P��c�=%�D4~hqi�}L��!i�{�Q�6�@�b3egmDi0�KO����4��a���������YM}���C+u ���]@�,�ɣ.����h��ۨ�>���7�m</�O�ܞ��c+u8��:M���[=��--�/��6�,x�(KKw�Uٷ�e�N��o9Q���R\����s�q�Ie�G��ǉ�7q�W�X�	jW�h4�c��o���G������ ()0%Fș�s'�GЯ��'BaՇ�6I����3��c���ȟ#W�\�/3�M1��Ͷ2��܈_� ��wOg�op�40=��q�r�2�\�.���z��B�cj0��\v��QC��7?�0ִ�3�'8�Y�q���_l�-��,�Ś�aN�_%A����ٽO#u��#z5p+ ��I�׭=W�8&� 50=���[Q}�����YV�.�����V�f?��M��piޱ��0���#��%��b>kI6��6>B��q��fOڕ{4�T��R�AX��@��-��|x�{�ѝ�e(�#�9%�t�Ǧ�ߊ�� ��OF�(D�*�ߐ̦F˸I��1n9H.�;�1x]���Isp*v 6+��	�h�wz�{���3�7��秤���Jy�G��
�s��B~9��A$9�w�R4��jn��nb�xC�vI��H�3Nd����%�v��NU���@��H�Խ`�y��m�T�f�V�[!�K�ب �՞bY}��E�$��q���γ݇;%�,Mt�ﭠnX
[�y��B,_�����J1B��p�|U�яϒ�2�U��Py>�/��_�)��9_�B}��<V�\�5�-�bQ� i됶��:�AV���d�F�Vj������>	�F�A��SP`��<D����$ш��|�zM���;�BjWv�e�F+D�sZ�[ �
��.v��Q�$/�K��M��
�U����*)����r��oX�$��N���US~�h�P��{lWX�`�!�D��Q�p���ǫdw(��vw;?�)�~$yͭ*&A�QROQ0 *�D�w1��e�����>kMwь������-WJ"�FT]��
���o�C��-p� ;�z@�0�(�vƕ��u)B�ҧ(4�t���i)��m�O�4�X��%qp��3G�+J�!p!�U�28�%�������Lxk�9��O��Wu ���F���h!f�g�uw
I7�iF�p�3��$3�$�ذ�)�g@Y %���&�ջ�bf*�����{X�p��@�E�L@
����<8}����@�X����nu�{B��|��ړ��l݃I����^�\�|p��O1����||^�1J�>��`�R��p��(t<8D0��?��b���ʈ~Z����~�U�����=�jDn+���A�+ϣ��D$������A��)�W�xk�xel9@5��� �i�(pMA['��$�A�*�A�}]�3Zw�$ei�H���u�8���֚���4�̓��>5o��n(��)P�3��-4�+��� �ek;"��e�8z�,}T({�vӘ������G�*���$��um ��J�ٛ�>�l��wG)��mg��x;�����r]@��7��U� ��Q�.v mT6���j�j�RK׍���8H�t�-��AuS����7���l0�ǹ*줾��k%��A��)8 {��q����U*P�����o©����)l�����St&$ֻ��|
r�Ć��D�����W\�T�2:�d6�{I�s����"��c��;��L-��42���F��b>���O�_lY �P���D�Z�KQ���/b�l#��s �"!4_�\���:x��FW�/�¨���^w>J��H��g��(��HVL�e��O�؀^Iap��><]K
>���1�i�neF��,H3w0h:?�Y��e�oo��#=
�E�'gr�<�7�%�N%;�F��f����<�,vb�R"��tN�ڹ�"=��X'}�Q��{>�+Xt`W��0�G�������hٗ�'���h���ձ��Bآ�%M�������,T�:G�e��h�"����ɕьe�O���K��QE�,�.�Q���������x���0
�3��]�J��
QocJ��'�!��N���S�	��#�?�yY����Q�����@#��]�ǝ�r��9�t{�u��o�ij�ަ/$��F�ݼ��m���j��C��"��]  Q��;gO�z��z��5L,d:bq��^���C\ωL TU[N�T�+�Q���H�����P���y[����Fj�1%�Ba_��I�;����шu��Y��j�WI����H�ц���o���D$a:w��Y���R�ě`ߒbV����b�<�~L��Ӡ�U1��CR�</M;�@��~�]�b��G�"_{|H,p�|E6I���b�/0֝z.�Zd�����I	~�?_��P����Ƒ\�d��:���@۸�Gf���|����Ȗ��d�M��8<-�A����8*(��w &⸙[��WVi��эO�����[;.�n�p��+;G':�~������%��i�����t��k���߯ovf	��8��,�,��W�,�����@9��1���x��7��2��8n���z�ZO
_���pLT�lTΗh]����u�dR`�=�����q����Lq�$�q��aM뎶�<�Es�D�,��S�M e��[���o>s���,Uy[��_	�$����6�E���CB�\���P�K($�&"�i��E�!*��$�4L�����M%[��5w���6��M�g�Տ��}Q��a8`�gՌ��I`꙼���^�ؐ��*ɍu�G�i�4�c=�)�m�FE�0&�>�p)�8��)�Z�,^�N���d:YUO�}�2d=%�I�d���0�
=�;�0Z��X�j��K��Œ�Q��h��� �����{8��kl�~��0�� ���H2��F���{h!�K�d�%��b�����՞�u�Tӳp����T?�Q��)�F���p~���g"v���[�#��{a�Y��j
�I��m�d/d{SL�5�t����,S	�C;Yx���ő߻l��@:�%�,]�=�7W�f>�@[�˥kysp��M�s�7x�v��6��}�=èg�)�qh���ODBTP���N�U`���`P���⬂���\ߣSAX>|�)�UDӰ���P�͐Ns}���őtI]Yłs�q�jB��p���P�T��^Q�oި�&�5Q���N�(����K�-T#U�h�}��/m8R^{dH�����i0��	����%���C�$����)
&�
,�������=��9K ��編\>(?/	��=A��k�'�e�J֍c0V0�ԩ��%G|��D�GD}�^��Sl��oU$~Q8S�)C �ӆ`R��qO.T�ay�3�:�xW	|.� ��:�˴��x��M�Ɨ��ݠ�����b3�M�j3�;-��3=�Y	�^����W�a�S�R��=3e˜���y�a5�3I����˶�Ƨ�����ha��^����N��r-G�� j�[���ux��M$C^A�3g1�_�s���
?b �@y���æ�E�-w�c�'��϶|���ʐ
`���ȟX'�b�!Tg4����=S�X�RO�B4�2�W�W;��zx���l�o5��ܿ��bv�`��'��xA���)	�I��,�~�,�޸(� �}� ��C����~���>�����$��QY��S�~51�?�	��J�<�6%j�T`�rF�������`��ظ���M�DÎ��F��.���G�S���0Q2oeX�)*�;b�K�V��ܽ٤�����R�+��:��\x�-���,�#e~8s2���ni�v�<$�B��
ЃZ��p(:�o���]<�����V���[L�u���z�6�M�#���Gf���TK����K�`��6#�QH� ���U6&���: ��z�d<����� 6��H���80UI@�������9N��6�mB��	�ũ&�Y�0{��1���c�4�Kh��K�i���Ӟ���{ �o+����v6��b`��3|����J������4�ك�������
+��7��pH�j��D��M1�3kR�/���ֺ�]�q���<@�0ߌ�f8��`1��D	Ƹ���cd��ķ<��<uluJ�s��K���
�����b�D��\
NX뱂\�.�?J{�Q�`#]N)˚zFj䐬�fY`cP��aǯ�YkX�0�$��YS��GE�L�O�s�Hnm�>�纼	u��!�	� ���=�"o	�r��G���nl�⼌�Q)$��Bh��s.Sh'�!ncK~��	d;(߲i��ڲ�7W�)RL�М�b+��7`/�^�5�d�?��#j����D�m�;�*����R�]%���Π�L���O�p������a0ӣ߀�B���;��>���݄T���W���:�&�,��g�"�7(��p��aΦ��c��V���_�L�)!�>	ۨ��M��mc~�N��1nl��_����I�x�F	�	(C���PV�{�<��	Jc���z��jZJ:�B\RP�����J��+����n�M9M�d?a���{� А�kr�/�Rܚ�]#�W�0��>�E�O���<�9���\����-��f~����,�F�=[m�T��P�
%�f�ԎT�|�Lh��+����vY7��Y5D��5%1��2g�r��A��bJm���G���E���s�����|R�Z�u�F�����Mt�|��vV�_dI����d���XzJ��E��Fҵ��a,�;��O3�����|�@�z
��'�����&V�ɧZ}X�_�0<vF��q�>�\:�vذ�:V�l��  �qjy�%���I�#{��(���_ y��m)G����"7dZD�������=+�}�}O�{q_�$�������[�A�3'b�E���9@��I���;e?��齛3}=���=oW6~X�X����~�-NN^�r���?��+ea�_��V�?� ��%��.��
��P��)(��}�_���C(�E�l|/f�*���,��#��5EKN�,V)a� �(�E��5[�<����I�,h��6�T��g|��v$�H����t&�=�#I��*K��Ȋ��b;�}wL�q�W��Z�_E�,N�����i���|P�T��0H �SW��c�`���5 &j���^a��
���0�������#	��(Q��N��2�n"��+S�@d��Un@4����4-��;\�B;�h�֋^���o��%��ѯZ&G��-<�F�j�M��Q����N��P>qY����)Ǻs�w�P4�Gd�Y���v��Q�y,�}%K2{5gsd�R��ϟ�� o�K�b2����1�`<����S�x2��TL<��J����z�o�`������h��P9m����>e�]��D��̕��V�/�k�颾�H��s	������W�;a�^"�U�6"Jр�EIy.���Fj`����_�꺜�7�ؓ��l(M�Щ�������=ˈ���#̝p�a�]�����{He��}I=�V,�Ģ�-R��&��N$6K����NF��(�w�R	���4��_K�Q�؏���!��"BPv�lp��ʙS��eѵ��+8g�N���L%���\*>"� L �Y#l��Ԧ��v���;@��8\�8��zO����=(X6?�� �E��ogz�w��Ѐ9��?a�B��r��#�"�����|�G�&��U�7A|���_@0 $_0V�X�%����������bI�}?O�6��pҘb�٪}$�b܈�� Y��H��!�D&"l�-����ʛu��_f_��X��U�LC�����xR6 ��Cj�����d��?�3�'Y�8M�CB�۳�NOt~�8#%�������\��L���e�v��G�C�|.lq�������Gl^�����m*u��qYZ'�8,��M Tp�YJݻ��Ŏ�PI�C�:�S�}�B�rS�
���@:*J�9x۹^v�*ek'���nRԯt���^	�BAe�z��kC�Ďn�*�rL�������A��K���gsN�%S��u��"��,G�uϒ5�`g�O^��{娵&e��Z7�X��b��Jv�-�.�F��!���qr_K����$f��O��Q��J
b��쿫3Π]yq�O<�2o�>VޏdXP�P���8�T����S �!?Zf"���!r��j��,��=o�O�E�u�(Tύ�Adi�x�����&�?�&t˔cZ����ƅ���̍��t��Y��ݧ��x%��(2�W�G����u�L:��������o����`�L]���޶����$:�LA`��q��$Yy����_�R$U�Z4���7N%��r�m�,9?AR�Y���cqH�C�0 ��^�$+� h�A������>���ό'�2�2*ʝ��@����M��H�s	E[ߏS�/�՝('�%��?�'�������'N0��%R鎈XZVB��c6��ި���I���L:����h�	�[��s��#d3�tx]<Q�����-��n�_l�Y�<7�·Tk�Y� ʷ-A��غo��/#拏m5�Ŏ�e|��&
��!g�F |�N�A��~Wlu	DkƟt��x�
�]c�$7�@��i�|p|�y��-����f��C.D�G�gaw�����7>ܠ�(���{��,�����R�E-zy=�h>Q՘���pÍc:�)�����V��QH,�˯��_�_2bi�Ld�-oa�u��.\fԊ�����zi���x�X6a�g�R�����O�4 ������u��zɜ����m4t�(���=��dzH��8)�4Q">'��'�'k�L) x�>�Ň�:.�$��hU�#.��1�A�\O��Zޖt�¦�I�VF�B'[G]8�F���OP��`������K�gV�(��ug{����+��Ӿ��@/�V��R�k��rvGa&���6G�r�'�"J�O�'��x5�8��%[���&�-{<z9�G$�1ѕ�Џݏ�\D�0�B)�r�-������N�G�a���F�{�+а��V2�&�9a����a�� ۀ�,�Z_ҩ/�P�p?\���w3i+��Ӕ[���T��� �:N�I��k�~�d�I�F ��ܡpcYr�1��6p�tPq�B��V�(��XR0&�<�X.��E�l�����/���8a3���vC���xBAS _^5u�����g饐v�W�������{�U���,Ȗ���C��������P[�7��eD<�2`!'v�
{Pf�7�y�~u���<�#ſd��Z<����^*���8.�VjD8�)]�Z���[�KC|�5�A�^whQ:��mg}G��th����v؃��9_���"�Y���zt�,	��Y�o.�-�Xr� ��lp���\��-u8��z�t%�oI�㤊M �#��}��l���*�,	mm`����f䖝n\v��ͣ��d>	�B�d��lA��h�ߎ}bz�����{��� z*|?�j�T�����f\�"\��FOI\;Dd(�y6�wp�r�y�+�W��T�D ��Y�K#P�c���1a �݅�R�G��|��Hv���{W�4��(�*ꅇ����;����`^��t%#���jh� ��@�Ӻ W��j�BG�"~ �4�xJ�@��^vr#��zF_��g�wt�#��5<����:��&�!��O֚U������@�Wg�_�X��*�kQ��"������}�ͩB�g�3p{�/<��[�����q�85�K����T8Zs>깖�iQ��HO�h����)�q*`~҇q@1�4�&q��ܾ�mj�,Í>�iqt����1�V���I ����l�XOj�}J�d���� �����f����FF�=���i9w[/��Z��<(����&=�}��y7��,�Q�����8��� =�f��+@ƻ��|��%w���w��J�S�%q>zL<�Ί�H�X�h�ƎZ'Կz�p�,�K{��=1��Uom�o�\΋w�!�v��S�6=V dc�;��i#�������i�T!>,V���@ҏ�sQv�5�-� m���r{@r,&� O���2,�~������� ژ� s	ȋ(��8X�K�N�*�[�H���}BIB�q�uE9V����-M�剦^t�~K�Y���#G�c�ŝ�����c���oi�e�E��a��{KH����x�=؍�WI���aT|x�RG$���!�<M�5F��`�٤b�V�V��]��|�g��jL䎜��@�}�uNN;;�(鼭=��� u�ۆ$N S��-}�&"9E�p��G�d5�fR����y
��X$��V4Y��K��	�ʄmq�2�#���`{Z�f˹�&�*���2w�Z����f�t<��P�nb����m���(<����3���D�@:��-8�;�w&��c��!L*#�^u5Ͷ�'(`���l�]s�f�D�SK7�/�GG垖[{/BO��ْ���F��?8�>J)�3�~����/1D~}����Ujׁ2c���'�Y(5ap�����v�LD�j��ϯ�袙ax���nwZL��Qʃ_�A�a�YAu\�N���;��F�8}�HKP풬�w�IfS���=�U�-�����US��
�(�h����Z.����*N3�x�+��sW@��hP�Ư�q�G����	���vk��VW��T�;{kX &(Q>3(h�= ��h�,�!���@9�ֳhe* ��H���7�a������ǒ�$�~�x(@���`JF����K[�rw���pPF�J�r�癛�4ph�//�Num�Z���Oe�P����E�F%ZQeq~��"龁��;�t)�sY�(���zkh
�t�0N�eA�LXF�,��;U�3�/? o��d8b6�L&�x]#c�9[˵
	�h�ml]O�$�;���E[j��]�?~�,%�T�i�X���J,7.�c"h6ã�wAa��aHg�F]�+}t6w'��.�/���yϋ�C���� !��}�v6@~�C+sBv��A�D2.�W�3�O��̜eί_���m;��cXY�rJ
�Ur(�8�����1�/��W��3����bf���w�N:	~�(�|����"��D�$0�T��84��T1y�1u�g����a���� q�o��]�i�{�To-�����R�DRў���I���?{~��P	AlP
<2e:��1�⋾$ ��l&����c����ܪ�^gK�w�0�Ίa�?>TF3�2o�k���������vض-����uˉ���ğ`�[*�4sځ�<q��N��� U���'k��Neޝ�"�4~�����2_Ջ��-��:�,�C��廟�"F ]F`�H�e��I��E�s��Lʎ��OE S>R.Éx�z8 �S?I��U(��7���!������5W4�.����n�!k�s�m����\-�d�ת�4�a�$���|�u�:]JXNv�BbX϶a��^؛����o���^D�n��Yxz��!V�*- �<>��k;�:4�|_�&���4��,q�H(������VW �`_���Q蚳�1O�x�AV�b1�ߊ�b��*���ڵw��@��y����t��SȰnZ��-��#�
��|�,�Ud{�V�se���Ba���S��1����iP^�(+�QS��H&%I��Y�sG�=*��;�I�������vMڝ�5r���#̡ �K����)�X."�.ӏe�_�n��nǵ���X�O�������:�l
:صs{� {�	�{_[��pt+<�Į�
'ۅ�稯R��2�\���N���wsW�d�@�q?W�!$�H2������0�2��|�_���d�DٓrS�h"x(��X|�$���@�p����Գ�!B�O�Z�=�d��mb���}�z��b�t��f!�G���Y1T N�X��~}�Qz*]�it:?�WK��>5���R��ɯ���W�dodxm�����Zގ/�#�Q0(��G�}�2/��k��B�A���A�P8������yD|Pw���>H�< ��b
b��S��d�q���Bl��%�r<L�7�v�౤s������82{��Ȭ����]����5��:�C��Nw�v�cH$,���@k� ���#����wN*$�P�x��;�jr�L�.VZ�tZa�S��(� �_�/�y�^����ݖ(n ��u~�"u������.�����|�[y�<8dV�	��S�5����Z��(
�f�I��.�^N���)�H�|W�R�-%��i&֋?H"�n|4�œ�R%W��(�flyͮR��'Q�&b�.jk�
_J̩%����G�bi�I܍�=��Y�3������5��(s~�'0�[g�;�f8'�/���ж��8�Y��>��Wq۔Ɍќb#-rg����{k����*��am{�&�穟}��h{L.��Xο���?y
ko�^�$�G���^�,��zn�}�>��)���ц�:C��ܟ�KrDq_��|$�Ɣ�S�<?HU����hխ���̻1��e���GSW0F�q!�:�6��Ҟ�B��dp?'��:aNt��xb��1!��c��a��Z�qy�%\ą6 S&�M��k�-.m�$�k�I�:��|�����g�	?)����e��["`7OHǽ�j�����������΅">	��
�?O�|�\ˎ�{�K�9���)�+�jq����ce����>�u@��y��}	�A<�B�s����?c�i�+D*��F�s�����B�]�]�炃:��"��|0��6Q1��Y%s� XE�j����i'���I;]y+'��M��i��D2�.s����;J��^�h��f}+̴�QV&�@N9����t9١���S�GM��@fq�u}{���X_����S������c��8Եف&?>8�j�����Ո�PiQ�i���ATv�*8�t�M�ssg��[!(��D�I/0E���%_��+���������tEd4a�,u7c��	������V�l�J���z�h>#�춇{�:@��| i��Ѣ4 Y�|)��7�ɺ��W[���{�1}�I	�e�����ey��b8�'m�s#٨�����컨�{��ɩ�:{BFoa9Vn(ti��8rH:�R��mZ���t}�T�3_��	 Ǌ~7ӝ:g�ǋ�S[BϜs׽��*<�N��ܚX��g�cb�$���k�0��[/	����Z�=�<o�H�ZZm�:�--�]�*K"���� �:�Ù4���Sr�_�&��c�r�h�0�z5��l�|��Z��Hq�qx?�{.��{uhs���Ff\��W\�%;-�T�<-/�J��q�^`����鿿����ͱ�!C�YuJ�ZT����ƶ�Ő����`�F�ɨ�����Nܒ�
�#�>����<hm~��%M���!+�
��헝O�8����?�wn÷g�����:��C\�՘�X*�9+#��P���nr�,ӯ�	7
���apv�%�l�%�[�5���ͫc���l�`-��������׺t�
з/%��܀s����3��I�bX�w	�	��V������|T�=]9�'�0���b�V�%�������m�jU(�Lp�J=o���.�&rO�P^_3(����C��2Z0A��l�IPK'I5T��w|7� �;-U��2�u0j�8����������"�?�C�̑��L�ubҗȹ<�R����nL*xRlV/��\+�<����`����Qq��!�˚��߼=�����B�*W��/������Fw	�F�!�!��Zޏ�g���H�^��ߨۿ��o�']<}9#ze-����f����(F���6>ɼ�ޅԚ58��J�\p^�Ń��aF�?����v�~��AZ��vn�j�,Z=�z���\�P&����z'�N}�Zb�����F*/�Y̱�Ôb �X��!HvB���e|٩�@W��m8�[�{B��<��=�4��?.Yۖ1����WM���1�ʭ�8SaB5���=d���.0-�gX������cS���p��p���R���֤(#M��	����@x��@�/,
4�uC��AAo��l� u�kƯ���J���܀�>��$�ZWX���/�=X�֋+�pv�`�ٜ䵆%�P3޿ga�ܠ������J=���N�˰�V�Ș�Z~M�9Jf!��4lY�?r�~	Dr��˸X����Ѳ棑���	.�@���]k�R�%-�-Y��g|���k���F���'?�����w�����wI�䨚���d���i��(}����QЊ������v�q�_���㝆��C� �����w>��&VV��啫�hC�V���'�L$���?��?�@_��$�"K�7��:R�m�R�#T�Q�������+v�
k�u���J�����U*]�����ӡ(�8��@�	:�Ff�q5^..�"�|�س�m;���R�5S�t�f�W
X���!����5�!�3�t|u�tے�H��/�Ԙ�j��7����b-�!���q�uH��������+	���y>�
�L�_G��Ϊy�(7�&��k���	r݆~�������9��s�o_A#M��o����7�\���iL��E�7]�0�.z��1����;��zV���H��� Q2�_r�G�.@۬%sܲ*>��5w]ݳ*3�S6��t=Y�#��X�-�xm[�Z��i��qP����/��'��H�$�k�,"Er��K��.�Mw�������i�.��T�T�P�8�<��j���.-;d�=��#Qsy�/��F�ktf0?���(���v]����N7:������UG��  Z�a�#����Ћ@E�i�%rw��r���(�3�-w}4,U]���e�湝,-O�єD���u3��7��m�>�Òד��vR�ϝ0?8�"e���)-Wu?�6u��O�kK=������s�j���ƀ���N@�Ǥ��7��N>�Q-��qz��mZ���ۧ�4RZ��Z��t�)�@˔29\8�[�Z��҃�틾!^�w����J=n�6hw�b>�}�G6��2�V��X�O�M�,�_Qk9��;�F��v`h\W*tE����Fg��NF�y�@v��������b��¾�G_�5�W�V�:��`�Z|B)J"J���LgD������Ҩ�"��H�K�S�<h�����آ$5߫�
۩/+��
�y�����	�$'F]s�Q���Ѝ���'_��G��aO��(���t�EBi�I@sA�|W."�����Q�\����y,I  Y��=����||s�78�Ƌ�#z�n����*
$���J$�=��I{�A��j^�c"���$�@�� ����vg4;+6��^6�\0p?��7��͏�w#!^�z����-��f2���B�NWr3�l:k�8�X�Ӓ�*�� n��,����S�h��Y������ʥ������ۢnEz���$�H�3X�cO��;�eY(��%+K���8ڻ��f��tϱ�'���HW��D��1�95� ��.^�j���|/^�Ve�Q��#�7)M�*mR���(A�Wg�`�-��C?���脺Z�Rvp���b���7�S�h5�-[�i`�����My�{3��r�Z�FN���c�$%��a]�m��~����w��2f������	Ү����g�\����,a�h^F����5���"�����?Հܻ������
&�Vò+��z�0�(r�����_N�Ы�����X��Eb���*��F!Ҝb�$M���J�K5wܫKؙZ����~�[�D`�4��AX���u�eP��s��_s����cL�PC&�1WN�US�^]����?��ɽFy�!�gq�#�x5Xl��,U"w��p���z4
e	� L�*}�[�z�ѽ̆�.��2�o�Ɨ��%��ƿ�B��Ԥ,:�4�Y~�?S��w� A��N���g��"��T7OC0� �����G��*��XU8��bR��4��tbX�"Y
��Vp���i�"�G�NΨ�lS\���[Vh �,<�8W��x2Wa-R��@�:��!���PLV���7� oҢ�[�W������f�>P>
�[,����Vb�'��^T\���V?���w�x��0L�YW�WS�Dk�#�J�!��4�4.�	bͽu��
T�B/:��n�"ɨ3$
1I��J�H��v�u{�I=�)��;�7��ݫ�T��G0a�E8)?�_Q^����>7x���9��萁΂=�2�Ͼ0���!�Uj�ɦ%(06Y|��T�s���T�a��` I��l;O�Oxm�/����A�<v)nZ�������$��?�^?~�􏩐��2^Ǯc�p�<�O�����{j�.��F�7hh��[�˫�|˵�����濠�%���Fޘ}.��;�S��q�YH
;#l�CޮT���I�9w���P�&*I)߅N���c�4��gH��+�57C���0꠱X���|�����N��5�L�8v���t%�����Ï�4���A)	m���A�Y1���q���}#��nQp�S�M�
�F�(�[+���ecWlLq=��cH�ia�B����e�T�:E�����f!��,6�0�Zp���m ;�6�=�A	+��E��Z�~XTlDx;� �9���wd�Ȫu��QM���?���m�B�g���r�H+V�Q���ڬ�0јg-���{�>�jfȢ� ;UG���2�֢���4emd�9��q��/ų`�(��J6�EQQo�}MQ8��-���3r����u��2���)��W�or�����$!V��M2��Lf7��@�+��A7!!.�Q����� -�&� ��N�J���:��$�����5{��/%	�yt����o�:PC<n�k�f�Z"���X$J�����{xib�Rh��<w��<]�	�U�չ��9r��.ڍ� �a/�����ka`�,�cf�b�A` i�B�7q�ܵy��q��ՄO�����mrS���_�Ʈ��CJ���ȌZ˶�&�!�fq>݃�<��������<��7�}U�?�U�f�S�J�B�b7/��G1��Mܑ6�"ie�w$r�:7� p��Q��}�s��!,����3߮��t�I鿱9)�Fl�~{�Zo�^���;���@(�*�_ꦤ���;�`���=��7���<�O�'T��> @ �{FA⒋gg_��O�w���S����_/\�"�X�kb�x�������I���ap�/wM�]"��m'�s��z��y��f�tIi��0�}�y���j�����S���_fΑTᒩ�L� �V̓&LC�a�B\j�>������B�tҹ��ٯ��g�%�*��2È7BF�q��� 60�(iV�{P>��4F�GwG�5v�q��?2��eлbۓ.,z��C�&���ʙ�C��u����"Z9�����`���'~b)�7X�O^�̨� �!���3$�B)i�οQ��z$ǫfg8D�N�Kt2\΅_B�׉̓���) N8?��U���+������7)'�갥?���h�	�����3��Ր�(����sB&��u���� s?D�s�A�$-��:�G�Ÿp��Ǡ��b�A��š����E���%b�1�|�� U������0�l��sخ>`��Xt��eڀā������qX*�<i�MӁ����,��S�^�yw>1�3��{x|c�$cU�����c	u��_p�T�#Eju��`�|�5y0m=�]��͞�A�s��t�����us��-�m�&h�a����ף�k��(ީ��j�+�nd�ƖJ=&�_�\/����0$3 ��ch�Pc�q ��/�T�3Luਠ���{t[�a��Έ�mٺ�V�67$Mt��`pZz�*�Dյ�οI9_� e���]N+c����ǩz�\��09���!/R �m=�Ɓ6ڦO$�X����i8��K�ب�0�	%��l+ ���;���9@�;�Vp�4{D��_;O㩗���^8�����8����߾���_9�w��)�d���C���a��|�4Y�/�f���}�d`��]v�H9�������ҡ,���e������TT�9�A���˨)��1{I��o�I���.���yN*�֎�_A��w5��������"�G�/��XpFO��:�¼8}ꪹ�G����ֵC. +��S�EO�yr��F��E[�ԹNY�{�l����M����6`C;x�y�)x0`����(^4���Y י�Wo�����\�&�5�h���ׇ��#�I���Y�A;W�0 �;��%+G&��{�Z�&;��w���?, W1[}�$����08��j0�X�R�ߥΨb��l�t�V�[D��2���@�6@3��b[�$]��PG���l�./i�+�����n�2��N��$�2�I�J�^�"����)��ń6x���Hka+�5H���_KCx���+]����ÔĶD��D�\��ie�����xgp��(#��d+�jX}��p���c���s�zq�:�Mm��m�0]k��zݪ�t��b��HM�.~��o&�0{��b2�)1>R|����p����_����҅6�Zbk�цW��4�덦e��Z�� F�4\���P��3���7uo�,Bq�6���sj�� �9zf��x�h���3�����Xj6\��7R˦���C]D]���ܻ�Aj|��^��~Q<)����󤑤��1n�� Ľ��ۨ�aj8�U�s��g�"����v�0�c�~��-"V.n��8n
�`��"�GC���M�W�;�EZl�_�߭eu��eӞ�c����P��������m! }�X�T䒩Љ�`�_h�Ӥ-���x�w3�g3���Xv���L��\!�]��%�������i�.�rn��#a�Ms��������3ͪm]�t���F��QeV�4�*eTj��1<�'�%�LB���ޙ���3�Q;)����4����݁����`9����A��4�$��q|f?�S_4������^�����/P�*����Ȱ��KAS�2Ds�	OX�޹�"��,©RV��);5�F̨�[���{&����s>��Q)�0ߨm��{�LWd��A�q����Z�]��1�'	}�c�C*X�nζs}"���ѡ��Q֐k"?��,��{�]^-Go�f���r¾�� .�������O+H��܊��T��xƗ�l���[3aRӐ%�L[�
M�r����e=��]ڍ�.�v�54���x����q�A�3����yJ������b���W�0ݯ@ ��ˁ���<Ȧ8�U�$=5�zu�<�����a8>���0�r�5V�ܠ�@�8��n����CT�e��"�v	�J0�V����ZI��aw�l@	��Nj}@J�z���Rk?FKT��q���J�X�$��a��%P�h�'$��l�q�Z�+�7�jY���y�f8jOI�a�4��FR���}�յ��3����w"|�C�n+b~ӛ��ZÑh̨�������P���l�Vfk�X݆l%V���c�kN�X�/ޫh)QDF��}ȍ�LFi2G�iCnv=,�����*#Y�7�PC�y)z���s���Х����T��ء�*Œ��{W�f�~w<',���`YF��ju�y�����`&$T�ѹ�s�_�����T▗^?�Z0,��F:�c�C,�&F��,��A�K��ı���&ټZF�z���w"�l�m;��I!�BK2�%��vj?YnP;n ���5��L��e��(
�)�m�}$j�^cN��s莰s����,�b*��a�z��q�����׺8�<�mzH��(�3�c
Mr�r0X�cZ7�Ҽ4�T�o�k���6���~�e[r[(��hB��3����e��K�%�!�te0��54�}Y�N��Vx��/3�ŵ7S^?��Jo����UF��5�Y]��s8T1��2�VĊ*"Fc�� mƬM;i��NN���Cw������N��W�[p���;�=�+�Z�D*M���d`�q�O5��X����	��&��\wպy�Խ{[�4�
w��.U������1;������4�!s����(u�37t�	<�K��QB��M6�j�`8���Ɇu��t����}�]e@-�5�@�4���A�\-l�61n��H��R�(}k�����{���SϜ���_tj��LV\+��>V�k��E暏�YW_R4���[����_V@2�P�&k<�t�Y��=�p�e!�g��G+�.D� �-����@����߮e]���fY�Cߘ5|d��w-M��Ĳ����t��\�|�"��=����
�)�,�=��2�� �JdFM�������)�?��c���A��4sQ�.�r���n*���F�!4NT8yt�7����c��}�u��o֫�1ͥ#K~ؤ��_��#���HM��^��W�,w����k�rx�g�ن������Zp��x����/yZ�N��3)�~�	�	���NC�g�j����I��p3Ԋ�.ؽ�n�4��M�рqr��yɠ��vs� F_�N4�z98��V�Ċ��Ge�3�!5R���[���@m;�CB�@17�N $x*f- �Z�~��5�)ނ�AF7AO㜸�'��iT���)c��e{�2Y��JD���  )q|�� G�b���Q��y,�;��{�a��5�����5cG^���{�E��w��_�䲹����ˮ���^A�x>��4Ţ��?��)�W��z����?~\�8��d�ӥ��z�rç���3�yV��w���x�o5C���~g��lHC���������c�S
4|G���ֳ�i��;�s�O�x=e��4내�Y�e�?�r�C��$�U9���LR���q���nB�Q0�V|�8��2b ��lpn��	�(�fG`�� �$k%�ʅ��-��^���Ԯ������Z�ǃ���oJ*�L溦�ǚD�\��<��4B錯3#��ih@o�P�o�f�Iq�io3*F�p��d_�+H�I���D�/bY��^H�w��s2��1�۫�_�&�?]4�~�1 �
�mB_�O�}�?�����9�\�Y �ױg�=N�(��寜�q��v	���Cp�G��~�Ӧ��cT�Fx�xT)���u-�X�����Z<dC����Yz �>N�k����b��,� c�9Y-c���y��p�m0��	�Z�*`��W�\˙��������;�)���m��l�� ��r��GԵ��`΂��;�~D&*tgܧz��R��|�؍8���4�3�Fo0P �EE��cƻ�eKA�1���Tzҹ�����
f������N��0�������2����/(!�@jo� �"�'�g�Of�Xׯ��^`����)�sl�/��)�h*&L��|�M�����P�nvSB�Q$�r��T2�)���bRQ���:�Lo��=vnª-�<�M��Ws!���JN�6820y����o���C�8h��"*�'��Y�A q���S�@B�2�ZO}1�׼���w[�Z��
8>�u�4Ot�0�:�8�X�-���ך�������d��P%!��*y*H|s��/��?�}]��o�;�i��#�6�9���;��9�I�-9�h6�@�fh�l'deʊ���oq�$��Uږ��T�G��G̠B7E��hц6�n$WU+����t�ܩ1>
/+�^KF�w�D��@�����C�j�e\2S��=�8T�.pGpf�t.4�dp��P�1��@W$�7�,}���
q�K���r)��H.��fY.��Q���M�[
f�?':��PU�]{�)�W�Dd�g*����H��{���1W�o�Y�>:����r�Al�0>A�y1�����Kv��W=��(gg�-��V����N�Ο���ʒmqŰd!~L��K?�7��Z_���T�T���e�ݧ�܋7��^�.
D��w1	9���E�0�8�i����������}���]����ë�6��J���;�&��؞����j�����B&�z�S��r����F����[$�h[����|7�=TPΘ��E�\����뾭�*4%w����m������q!�o���(��[b�iJC"�`ZB�,����+؈.歰hL��Ü,��l$�DEf�Qe�5~���S��!���u�ek�-���	��o�� �(��x`kEٟf�l���|?U�;�� �4+���C�~�Us�O�k����ӂ_KUZ�Alذ�ڦ43R�3�`|����7����/Yݕ�A!�l�29$cRs��L�v��H� �#�=T��7e���\�����b��/j��t=�#�;�#��������7�qi(x$S��b�Ȋ'B���f@N?8����e�U�ޝ��b�K~��#���-t�0y6Vv���譖69͢ӆ�/Z���d����a�G�X��LL������n��F��o��v���t�o.0W�j�����l���MG��e�����_�v1m9�u��4�Z#�~&wv4"0	�%�]g��IŽV�qh�E4��lǅ��.������L&0,��?���C�_q{�8�M>�P���I��W��.���_��)�tU D��YG��\��5{B�YDh0�辎�~��8�H�|���ʤOPc?z~�K�\��I�F�"N��~Ў��M��7�'t�I~�t��	tt��M��׼�^]�9b��?�~�'h����Ԇ!1������[�;_��(jKC��n8��4l�W�a��[��>��&�g=#R`�9h��K���B�����[^�- �o�":ȄBH(:�̐�����o�L���.�%h�ӐKnN���u�I�=,�׳uW�y;�epWw-�z�34]��V�3>����_�����A`�b1���YV�6��R�T	�������� �+:w�7��P� /���'�Q}{��Uܖxn��Hm����OϷ\��`4_?�J�\S���x|U�̀��R>�R��C�Z��k�J�����K%�� 5Xs\����C߿��l0�"=YK�a#x��]�_�����
�[����ttx��H=��n�P m�]8�\nb�rYs`6=?]�6B�ԁV�g�M�ܺ�bb���K~��-h�g��D��+�:�o6dj�09�E�j�1멦g5�3Vu��p�bc�X������g�[ ���㦋�5�1�����l{�3���$��T]�<�(�Oeud�g�'4��䵡6�����=P/�}�Y���A�����c�KI�추��Sե.PHz Ǘ��c���ݿ�RV|���N�9Gn��Ƹ�L��:)�nH�Wt����� �S*��e� �[J�q0���1��F�u>��X&��g��Y�q.�5��pU%��6anV_�-D� O�<��b8qf,�)�#���d���҈����I��G���b�b4+��d쟹塗�����uLWZ���|>�!�����o�(���[J��<mxBP��w�̜&h ���r�fS	�h1�a65��� �j	�q����C�7�N��U��&j&���&{l��p{�Uz���3v��E�b�ZQ>��"D�@�.湃��n
i����>�$~Ύ�'�j�߷m�km^�ʲ ��~v2B�9�>[��s�ڪ�I�(�R9dT�֖ A2�o$��%�w4]�d�~,yy1N�w
�x�v��`�κt>�l���H	�}�?�lgË�z�k^ە��O��a��=���6> ��2�ҿ�s�j8���(|X�����P-����`�R�}���M9�5l���d��֪���"�1��.L��� �, �1��|��W��ȡ����hތ�) �,�È��;����x������1K_�VH�ʏš��XAR?hi���y?�sjB�_3�,G�����Ժ��HJ�ޙ�Z�B뺽��?x͇�-�4ɪH�N���,��ΦW���� >Gd��X�tUd�-�@QI\������R����=��o�}��<�{ٶ9j����TO����� w5/Pf�����pNPi/v�'���xW�L�L�����皰(�B#}����$*g!��c:d�>����� ~O0h2���_s�r]� Uf`���F� �QCB<��k�0|����;H�S��gO���[
i�Gs�@�4�&\M^��8��J{�h���LW�y&5&f�b��:������b�쥷�q�y��s+cе�"VE��\�{4 L4��H
3I���@���k�Q��~}m�K�h1C�9JQ�+�	�k�}[���V��d�3�ش1Z��ԃ2����r�j@r�uN�\1l�ifA��*�Nŭv�}9�S��G� �g=ţ#cIw���� ����gwH�:Xe�7�����J��4��NgF=TTo �Y���9��8}6��\e
Ytd,�Ι����a+s�� �/ ������g[.�[�VZ��Ԥ�'2�أ�M0�a�Zu'�_[ZC�c�`�X��5e�A�6Cx�(i!
����\��Lf�
*Z��BV�SqpU~!����^���?�[�J ��Ƴ���%.�˽͠���\��R�)��`�Һ��Py�.D��c���|�����7��%O��&�󂦑&�2U%�ߚ���_KMSצ�%t�@b�9�0O���-�7	�ʯjd�Y�J����'����>��(3��k�3���t>�V�[V��r"W��c����C�m0I%��s%�f�ʉOP��W��<�$�O��� ��4̡B�S�i�]Dt�������N(�b�Ҏp՞52,�ғMM��稔�u��^����Y���T�+%�_Rފ�U�]��r���EX��]+���!2���q�S��������9��n���&\?�D�fTB�VR��YG�A�����@4�N��!���b5�V����=X�oJi��[Ġ�Xw��B,�&��'�[ּ��P��g�Dq��#��C�K) nbtm�C�5�g�U晇O|"��U��b@�H'7i��赇fF$3qg>O�#{2��Z��[�WR�\���+�1+?���rJς���N�T�;ث	�t;2F0\��ŷPw�����~#�&6���c�y�d�ҤF|ѣco:�0Z"U{�c=�*Ϳ*��x��d�����������T�F�9_��`����P�9'�8�Å+Fj(�;��E5ݬ��M�+���,�О"�ҥ��:�O�aW���Ƶ��g5I��j���h��l��Q(���bۊ���Κ�@��ֻ���*���Z�m���<��db�S��'�Mx�Z3%�tk����q+d�簽x�q�PȺd�+��EZ�MJc�F�[S��)YL��k��x��	;kB͓ԦB_/U!+��)�-�'��s��(c'��=��[���%�vG��\G��e12�~#B'ÌD؛�}�W�z�i?����8�hAZ���59`0���[�	�����s����܀�u��F1���w����KnphRM�\��E���v����}<�Д��6�0�L���"�Q>W� 
whV쒤�R���t��9Ry�����R�1�o6�ߡ��N��K�0��u��V"���Dνv�S��Q���$^�i�U���e4cg��	|��*�?�{I���d�8J(�e�4�(2�ݼ��͵y���'�9.U�_L�k /���{�~��,䚰$��@!T;�&[l2��-6�j��W"��I�T|	N�Ju+j;���ƪ˭��5��T�PD��%Qa�$��&��{�ij��{4b�/���զ�ɏ
g���Z�H>ǀ^��W���-٦�ԏ٧�o�ՙ\Bcd�1�X �����R=���Ţ���W��}:�R�#uu�a
Ns�Y�ܹ�����uC!V!����)�Vܹ���P1oZ�{�4�O$@h����D�p����^y�O`p転*�"2�\c*�]�t�Ǯ�
!e�vcoo����-��\ƽ�jkxtl!t�NWC$<�{#MB%b",u|�8���7�x�|�h���a�_uB˕���X>��8@�?��4|��o�'�HQ<������ĥ������t����E���4�U��_�M^��t��9���c1aX�ŝ�df�,PjpC���'�.�[�\��I�C�o
��4��S�@��ݝ,��N"+;X��q�)f�L�ƠR9@���N��%�9��f^���c��S:G��OT�� ,@`�"M��*J�T��1��Sc�J,��<xA����'�ڱ2�3>M71B;����"�?�{�𓑚���{@�&fCxf�S9���v-��;�V
n	'�-����ϔ�2��T�1H��G�~�����X����>�&c���I~л�M�w&�8=B��6��p��i�{'5e�(�6u���K��.%T6k��eJ��3��Hoj�{?`)l��?��,��jL���5,��z}=�p^)b��S�wv�t�~%E�ݻ�;,B�Pӧ���s�GwY�U��	����MXs�a-Vr>���\�귽y�e�]j�sْ���J'�wr+	�D�.�R=E}qWS�z�D���#Z�G�����'���'� x-�~Щ����( p�=��C̒xf�D4l�+���QF�U�
O�y
�[��u���W��K,����T^[�����&D��;9��R�o=�h�v����`Ģ6��eR%�^�EA�չ�\��>��L��w'9���Dv{碃�pb�2���@�|&(�N�o��J���n8�m�[Ը�-�ۘ3�dȎ<K�+7,�y��r�����H4����K�k*���3���g5����/[��ds����{p�Җ����$@��3�x���wrL�Ǝ�4�hn��!�I5ZS���GCr�&���P�SI�Ƽs���!��a��/ ���ʰ�t?��m��>� ���e�O��7)c�?<;�c��q� 2]�b0��+n��cN�P9��$zR}�4l!h��:�ס�;t8���w_��0X9�M�<��i�����
#�+��<�-La�!�3Px����>��#�f���LKTƝ�x��51���.�͊H���x \'���t!�ғtFbϝ���J -�&{�#���Pڈ��l�(���	�V��@�.x5��w��ǡ��/A�6�f���4]zo.b����)̚A��o��x)#�V>28e��}�q*Cj�L������y�^��q��k������g,J[�kPҜ���Pr��+���#�1D��P�~��R��/��d7�@C+��q�8��O���&q}qqS[�`QG49Hwv�L�U�w����UU�/d4�
�F�M���u�"ꄯ-딚�D���У)��o~�e#�&�|���L|K�G}�;^O+�y7�{��pJc5lAu̾9�$��$l]�!݇��Ε�#�yy)�4J�j)�"~����f��a���m�|���^�Fp�Zp�T�'Nw
?��'��,B��_���؂�?�7}r�,*5���
Ǫܕl�Mo�v������@ZJ��iɔ��?rZ�X5J�}��_l�J�3F|�� X��F
X,�L�ER�A�3ko)=�4P���^��YzB�0oK�]�k��Mqv��(��w�:�W��^�5�����AB#%Y�1�`��s����M)1EY��/8�r�e���n��rC�] W,Qo����O1<�\����Π������S���fP�9���i/�JYL7U��ƨ�I�(��j�g.���Y��1?x�������'%<��_fg����pR���_r�q�a��ؕݿ����Z��N{e7�^�
��V%�/+����I)��}� ES��R���d}6+��l�Ăib��%J�ƻ!�[Ɨ��̛��w��b���g=�i���c�P�޷��6��Κ�$u�O\�t���LP$[��o��$4]z�m�� �w�`[�Ioa�H,26ٮ;ZV�s�:#�>7����-���޳��D��i���fă�1Jc���9�8���	�}���6ڋ� �#��Zh��﯋;=9�Lk��qF��E@+��E-~���?�o1&���`�6��r��*v������^��� ��;|���>m��4F1z���çE�W��| �%"��5�������g�Y�K������oD��u�C����~m��H�
�������Fvm>U��8=��2#�_�0mlnO�C��Q(0k�ޱ�7�;��`�q�s�T덛��M�{'9�]�� ��WH���ǬzI�EmD1�/S�Fm���L�������S�?w~\�ŗ�N���ucѢ���x_��5W*��1�ݜ�H���\��a�1�Y�H��}�U��p%	<�nE<@)���e����n|�q������7��/W�z��c�Y�SD�`��|�:��i��^\�k�����m���B�v9	�ʭ(&F��G���<��~+��3��f�%�s'_]� !�	�^=A)���O�vQ�������zL����c�v�K��b�A�ٿ+��-����KѨ�Q�a�����Fr;����5�h�a�v������O2�38&7M��5�g�Q��2�\���¹�Kq���
$�Q\�ȁ8�1��L,sRq��I��;�?����,FF��t<��㹰ZyD�f�\��d��d)K0���sV����^���Ea�p3���U�	}>yt�M����οԑ��G�Z��V��/��&6�7V����^��V�S[�֥�c�k�j�M0���l�����	��}�4!z�Z$���U��61ѹ�q�@��z��~ pt��˂��1�e��(?V�:�XE�)�xt����Ť7��c���l˛��&{Ki!������Gr��s�IK}��&����(/GD˩C�J���tn����9�E��)0���8����x�z�z+4=����i̐].uV�Wr�h%��@._�M*=���D��,�1�~���W�§no�H�]�=eR�~�b��3��]�m�m�Ie	@�!aC������3��K���3ٞ׍9�����x��Q��)�Y� ��c�����ϥaO�h�F�"���
��(������%`��x_d��+�����`e
x0�7!�<e�I*��4(�}6�T�.9GIU|�z}�[Qi���
�؅ߦp1��?xv�R��ש���qF�;}�݇�ٷE)�!֕-�(�V�S7��o�U�g`��t�)�}���D/�y6+�Ll۟T7��+F��pI��Ѯ�
=����ݘ_��B@H:�W�h��[�~Hb0��(T�n�6�	0�{��Y��A�g7�C&��A���`�
���'i����w�{ME���T�T�%�ˈ��MzW�F^�>��)��y��P��h!����=|��� �ꕃ^�h���LaУw;Hl���U����@<����dRX��RA����po���E&��f-�$8����:��-���LI�/�u�a��p4|:�1��L�0����~�GL8���M���/r���	�c{f�]�zܩp�.>R����D��=5�X>]��"8LІvm^��ޅ��^|�ɮE���xcF�9}�}�t,y��G��Q�g�������@��*� ��~8G�����i�S~�~1Ւ��5�!�2+�$6�h����&�8��6X����#����z�k��:�a�'�����
T_�ҡ�:Ӥ;���Q���E�X�ǡ����_���_I �e���W��1UA����G
DF+&��r*Q'��3���bDd��}!��V2���nΊ4,������	$�%v.�K�U�_,s �N�����Xd&�ZK���^7�0�|k8f5�E'�ti��������z��u.�9:l̎E(dpJT@��wxE�F��������i/���#P�D�JU�R�R���'���n)��mo�ޫT�펑��v/qiӒFA�%�Y�����i���:j���〵#õu��O�h��r|�+��4ֽ�.��I�s�h�\���c.k�H���Cy��6H",T��Y�"w�����g�N�Z��>h_�@��J`R���Ĩ٪o?>��
�����m��T�i�/��0����6z�ě%���a#�a��L0��R�����S�r�Za���)���?T�<��OkҮꊻ���X�E��� ]�� �#^w��V�aJT��O��z1���%�w4S�k`SG����h%9�.�C��Q�_����Z4 ^Ů{���k�E���T����V�]�d����L���D>c��k��OQ)��v�����Lah�Ôx����K���}��2Y���nI� 1K����{�7���)G�Dڟɰ��=#сn�L�s�����e�F_C����Q�x4*J.�Ǽa�)��l�n֫��!r'6W1�/�|쥋 ��P��C*[�_8��zs�]c6T�퉯�x���r?��"�����Ly7	Z.����x���G|��T T���*	��p\MK���SJ�{h�|f��Q1����Y�k�t����Gu�x�lc`�贗֑��ӻ��?T���	�A͌J;O%o�*�xUTl� ��=�MO����	Ԇ�c�y8t���;�(?�5��_���Ǐ(������oJ�����2�����;���PP]_�H�]�t�L��H��/��h;��S�^{%&ֿ/�KY^R�X5�}��O&1i�V()��Ôԗ�f����@�/k���G UM� �{K-o��V�H��E�+y�T!vQ��C\�K�r�q����j2�/���!��P'�I|p�̓oa�t��?�ƷC	ώAτ��]��Z��r����x�CC�]j���Y�t��Z��B�7{��{Y?�q�e��-�>;���^�~��ܫpU����e�C�L�1�{ ��PoW�Z��tZ�������Ȱ�
|��Y��|��PQ������I���'4H���Ik��?����.o���Z�hV:�T���C����v��-J��3�}t��LDܧ6�ɒ8:��:Ba��-�R��f����'\j��ؘmv�J*}/��aW������~�/
��nH-Vz�X"7��Ңرt��WΖ\��^��MΝI��VWm�$�s���}�d������P���qX�?�+c�̢2�aM�I'�˿�����D�8Cۨ��r��
����GY\h�X9̀5qB]���u���?t���Yߊ�����g��kX���/�o)[Δ-ϸ�k�l7����hg��=ԙ �ek�A�(A@���yN�0�,�p� ���r�;�)�dМ���k�|,�)�i�n*|�{�����P*7U���5��b�t{+��qĉm������$��DJ/�$��/���#��?���GIf(Bq�Nǧ������8
���*��=M�?�(X�&���Dy�B����VN��E�v�^�ǲ<���cs�Em5Y�I��l=�vAz����-F&[������6�f,jmAOWR�P2���@�i��S���H2V�#.�H���h�γh�[�4���)���~����J ��~��?�����A��b�K�i�<�a�	��J}*X�VBImЌk�8��i�.�$kh��2 ����y�56��T���~��P>xfO"S��I�n	o��T����v�28k��� rֵ`���>����$���e�����?+O$ډ��'cM�SR
�6N�n�yu��f�k�vŰq�FP�WP�oh��݌d`+Tj�wK���1��E|ddq��k)�����
m��py{=�����&�(��iΦKУ�As����d#�NA��a��є�����d)���g�𣗐����5��m�FK�[�8Fw1?i�C
��_�Ֆ�0��x��y���7l��w�����0]f)t��<�����)p�g�����?5��k<��a��"Wj7��+�������#C���xz6E�r��z����U�q�%[SP"	��|J;P��n��A�$�vn��=ɫK��� T^ikÆ��F�����9���Q?4�咫�y͹�]+����)*-/����$�-�hɸ{�Y�#`��&"��[����������ɭ��] ��,fTx��9�\~%�2݀�����X�(v�V$���o�|�浀P�(-{�"T���� �����
�t�"�Uq��l&��� cZ?�H{�F�you.e��E��j��z9�b�9�?/ݴ�R���8kjd����e{�����Ո��F����"¦���k��g3�����
�a�+�cu_��tH�k/�
"��~�y[���E�t��9;jF�����.2c8�gЖ~����
fNE�*��ϥ�y8�f}2�z��>��.-df��*A���D2ҳo2p�����T�D�_��0�&�BQ�V�t�3��`�J���6&��u�-X�W�Հ���5R���2n	�%�.��Bp���ts̨K��3�&)��j���S*��a���.�5�vVH�]�J1(�R8����f�8A��Y���9A} 0�^�zP�$���Z5�M���?(�G2�t�צ�\H����W(x�f�vo�?0w��(w���y�Ӭ��٬):_��*M�gp)���6�]������rSTހqj �{��  ��9���G6arom?	}}��;C�$ͼTQ^��a�a���w%�(�u��8άB^���ط��W���P4hni��W���d�@RS��z���>�^@�� ��H�&�+�N �&WU�CD�*�Z;�:�)�F�T�u
~���D{�pOF!�l+�L����QyHE!�E>8XВ��VVÄ��^��T/ __ƙ�{�9�	ޡ8[?�0�"PiT��1G��m"��R��iwVR��U��<��1�yK��o`ɾ�Γ�#����)$�Pt�B��<˼m� 9����b<`����֖�MF0���� z�8.�!��ۗ��nڐ���َ9*�����S��ޥ�O=�fsA^��۵d�>AС�p���U�x����Q�2R�e&���f���2�W-�D//׋�m$-��k�I�6>�ѝ粰p�<�KÀ�<��gD1��W*N-"��)02��x�]�`��]ߩ���)�4AhM^���j�y�nd����5�~͈����q���ľKB� ������g���.�!��[�#O��|ǔX���k��6ku��CU.�4��AV��0�q_��Hq����p�A��Y�\ �.��.�e#�<9����ɻFR���>��#7�~���s���P�mBo���,��x��6�d�Y/,�0';9�!�b0�[{JbכG�	����?t��ш�>iRMy).�md3�Ks��u��b
��&+ܕ�s}̏_,�,�ʖ��2��Q��|�U��,Q9��aZc%
h�8�q�@��Ad|���.c����P�L90[|d�eo�HЩ�r(�uO*��3D0G�.L��$��i�ٙ�yVd���V���L��%΍*+m�T�0��w��V��[KΆOk��|ʾ!�sG��e5��9m�
�f�1r8�|3T��l�[�N<G8E] �\9|�o�����uf�;�?���cXe�e��M�
|�ˮ����Y����]���J���?�?B�D*k�u����n��*8��n�1,O7�P���$�����)N@A��T�~�8�[=�Y�O_oq?�j%ق{G��E�׻�yh.����0�(��	�N��g�[N�p�q���9�}����R{e>R�7B��P=˟ڿ�
�uh(�I-IY��/��2d��N�L9����0�o�G�ɕ��n�����,- ��ث���vY�ll�ȶv�EM�Nhd��,B6��m��
P���2|� �Ͷ��(Ɋ:�n�?�o�Eq�rR�]3#pk���f1��ũA��\�e7�/m�{�>�yW��$W�����v����b�Δ$@V��R�Ԟ��s�nCjf����đ8��s��FK��]q�̆;ܤ�ܩ�{�Q٣Ljf`��=�'��D�p��(/�ol@
�5�l	<�AW�5��P���{I��%�&�)�ni�t�A�*m���!֜uC�\�,�w�����U�.����ة�"���yĬ]o��Dr`�l��<.fr,�c��W2=���"��F���������YȻ~��s�q;暮�]�V#_D�0�ζ���٨����>�V� ������$?��ʹk���!n��"�c����FW���`*E�L�n��	�"���h��ۤ�
蹛�����k9���1<�wF���~�_̖�lZQ���ѶrA�&#�L�=�gxE�1i��z��[��20sV
�{?���=����F��4�w�\�m��es�r).�$}���-8�����zQFU9�V�y!�|�J.��Ŵ�Z<�w��NF����O��#ݭ/�;½uFn�`Y����O���[�z�S���}�P���1���-<dh5ŵ����E���b*���\���5��T�;v�BF]�&~�z�%&��%�ڄ��/����� � *f5�2"�"���2�.�����YٞLF��<��N�LBa��(��pI�AsR�(�8%�Y�U��[�D-�@�S�{2uYA�+�BqO(i�T#3OC��Fk�^��]ZLMS�0������b����3:��Y:�m��b�#$���)�j������e�Y�f��g�����U�[��Ŧ	���f�X�y�����{l�;e}�S�½C)���V9=A����%�|5�Z�!�~})�u�'�����;��X�� q�E2Ֆ�c��#���ʖ��p�rO��z=�K�e+S�.ë�MIPj��p@�)UBZLUf�:?o�*�����=z����\g���<Db��b˗"�3Z`Zc���i0��VB[t��ᐷ��i[M	�dv���r}�"2��1�#�G�2�!!��u~�o"V�S�h"�d��W�����˲;�L= �J�9!��Or֯�D�De�]M=�q��r:�$]X`Ki�����[ϡE��Eu��DSEC��v�?��p2�@j�4����X�����T���&ъ�{)��J#hh� �$p@5l����� ��"����Z5R?�+��Po;���,30	A'l�������
ZtZ�g��wn:�������/i���r�O�=RP��b�?�S2z��P<>���i b������M*ݴ��$ت�/�5�[|ˬ�1��X}q�=�F� ^���@'%��Y1-	c�`C���M��V�r]栧e�x^���L	ա���x'w?�/Xt��h���evq�����x�w��fI��.��ԓ�iڄ��_G��j3 ��MƂ�t������h��9>�[�F�<��C���ME�p$���������y�Z����ʁ�Iu����y;[���Lݮw=}�H�3`��/�t�r5����t����vE�-�4F��>�K���7%�o�F�`��1$����vT7u8��K6��0h��P�}Q�.�2�S��=�s@��Em�j��E�ΔrR���e������@�؉e1�2V������k���u�/r1T��+~�K�d	 ��h�`J�Ր��q��/�|�jZ��$~�*<@^�>���{�b#ag~���ǔve�}m�³�4#hXǗ*����Y��Q���H�P3h�{�QO˃kZ�I��a���
Ӕ���@0�e��x�$�^����yn�ض��@ \�U��l���iN��� Mu��W�������TZ0X�j��88� �,.#c����|�� ��_
�b��u�/S���a8T���3F6�@�	R����D��زS�(�E�(��_\'����]|��Q�r�SBh@��V��?�������^��0�˦�KGE�Qq�M�`�����2�S���A��t^�۰O%�|0�x+sž6���Zp��m�~�ݡ�$�6�����)ǥ'_�pź٣�%T6�9G9�:|w�G�ʏL���D��4H"v$�Ԯ��bǸ�%d��3o�rZޑ(��t���[�Р�(*A'D�ۖ�Ⲷ�N͖�:@���d����nq�/�Bci�z0w�	q��mT��|EG�������9���������yp�U�%��<��'��� ��v�7/L�1o�u;j)���b�Z�v�]7�� 2�~ ��Y���L�eZzMl��􊁰�.�bp�aJ� �H�^A@�@�\������cj�{��o���p�^g"lp\HC%��v4W����̛j)=��
1GW��\F� "hD�Y�V,į�F��U(=�C�,���zqoc45��uj�u���z���{>��S�d�����=	��B�_h�k��8@>?R= ��� ���b!U+�(����n��2˔�[*��R�+4�F����V��H�b�çU��*lA�q�VB,���x$�mC����|��h%ݫ�rs�^�%�8�{V~08є1��T|,jbv<#y(I���5�����߂�	�[ޣҀ>l{\��Sc혓؝���=�Q;���HA�f�"�آ����۹Y�?�_D=���[ܢ:�Wt�y��I�V'��bi�n�V�fG��؎�P(���5�-��$� ���	$�v���V���cA���Ь������J��t�〙�6ަ��`ٮ$�c*�E5 ��Q˸���o�̠�n@=�.�߂��x�6�`�r[����R��T�;^k���:d��%�����]X"N��O6>�[�"���Ě-�&C���$ptC%�(�ǋH<�C$�2�B�����b�P���ޠ^�ne���n�/���-
��6�St��"�6Gw���&ux#}$�y��)�nq��|$��qB�a͕ ˼�c$�u�vY���xvY��!�ͷ7��v�jd��=M�9���=���ݐ��b���N*jcj0��/�d9FlТ�ݖ$TΌ�sE=6/K��J�&"uT��J�0c��(����x�-VV�
�ײޔ�(��67H]m�g|-Bd��A�H3.7�U�y��44��l.�$�6����x�����4'��Rye�4���,�f�1�B�@�z"RoU�����ˇ��CӲ$��Y���h�@�__#��5Ag\?����(_5�-�oTi�D�/��d���XZ����	��9WN� �?GZ���r��՗�N&�s�����)J�rV�}�2�������#2-d�s�!��G3�Y��F�8}��:��A�?�6��YП*.��^��.pb��)H���} ^�#��H��~�$���i���®.l҈���,:V��4o-�E���j��b +�|qkC��ʘ��O� 	~��BA�z;/
�)]U���9�*��p�g�l��Y�%*Ȝw���� i���洐����~y�����-�7��=WòBmX���r�i'� {�a��
M4�%Ld,�;ԋ����1�n��?91�.l�!O^��j7�y�����`�r�ٟO��`w��*>��{�����A��FC������.Qܿ�s����(i�L7]��o�ɉMԠ��f��uQV�ɫ�pq2�����|�p}w�]�_�1�.�o�Ϩ4N6@¥l��J%�2��05)����d0�HքtACs��b�kCP0���ba�<߆�8Ӭ�m��ٵi��%5x�$�"�Т���bҁT���L\exs,����J�ez��蜤d�=m#�o��i8�ֿ�-�<�����B���}��+�g�U�	_I������#����gS�E�>O�:�!Kh��Cy�L����C���l��c�v��	����l�����E�� ��əGj�v�zɤ�;��[��7^K�b�p�V�2�';�nh[�@��f�w���7�1Sۉi�K$۔�p�w�cn�d �1�fǬ`t�E�U���h9<j�h��D֝���c���Ue@[��jY��*���r�9����[n�"�7��1���,�Ô6�9]�����{�>۳�l�Q�58ğC��� -�&������=�V\1	�1�3��^3O�o��1�p1o<3�i�{
�>���	�{��y�W�Od����ô84l#�R�)�kW�u�JofsZ+��a�{� ���[ƧvSn���蛣�q���V�E{��[
S^'�n.��+'\�W}��2k��G�wi^�~S�.OʮDq�X�ы��'~����Y�:'MJGgTƥ A���h^$����]$#UiK����}LZ��3�b��c��k����+� a�O� �"j���!z�vC�oQ*�O<?�&��2թ�d����
�6E]�̢b���"\�|��0�)�1&�P[�I���O��ڒ�i�Zʻ��w��0aMQ=����Qm����ee6�U�]�� �V�G���;�ml�����1��1��V�eM�-��wK�,F)«�&�x��G�ف�A�y!���3�vnJ�Hmz8ID���xRs�7ar��4Y㗱~�k�������5V
:O�@d��T�� �P	Í��U�EN���U�4	y���6��A���ѐF;��t�R�4.������F��v�p�~6so��c�� �W���L�C��9�h���u����MV�X�2ON��a*��SXE����'��V����G�K?t<\WۂZ��]ͭ��4��muΝ~~y�{��_���(=y�8�&J��&
�k����Fh8�ń�X�sJ���K:ĺh���C�ҧB)����yf�q��l q�v�I��F�J��&?�
�:}�KRD�sV�r���#.  �����4����B��c4�<R�n����!A�t"3��Ӧ��e%<_Y��P�@V7�o!a����bwNC����%ʶ����Ǧ��3�}�� �� u���>�Ȭ�ׄBv�V65\d�dg���/�Ak(�+�3 O��zp����!�H�?��ĺ�̛���gGO�Q������r����\�h����L�(�$Ğ|4p��1 7��:)N�$��N�G�K�xQ^{� ���M��ؕ�G߆B@
RV.���^��Iđ�)��ƶgG�e�eu��J$Ԍ r��>����Z�*�lӝvw[�
��Lq�8@<�#�J�3$\�"�õ����␶c8��q�,��)ڿ��2��Jyꇗ�� �����l:k<���1��!Qل��G�[����jx�.�ԡ��.b�q��j�x�93�BY�Sf���%/o������Fw�l��9��gG�Î2�B����E�gmG��l����D�^�iA	�����?����t��f���p��.��pЅF�MUv���C;uo�YV˘s2�0�=n���c���H�$�{e��qc�H[H|1��ІX��J���b�!A���N�t6��Iց2������b1Ϭ�ڄ�������2��V	�2�� ҁ��J����xr���B?�&%�?����XE�����0W��CNeT��TJ��F�Z�b''���3`���^e�A��T�o\�����\��jVy����`�}�g�|��'b8^ ���n�/t�H��
�X8���~��*A�]�7���$�x�׌����PSPP�+M��DZ
����ۜQ�^��nV}
	-^�		�����qa���]�"���]W�B��$ғ���|��t�O�r�o0m867�iA0��Va$`'�7����l>��&qZ����l��1��@"M�$~��0V}����y��.�/���y�����<�z���b�X����BBB;:<�=L��Jt��dw��f�RX�^a#�K�V�� �O��J+�[#1Y�y�AM�T�iF�H�w�f�O�>=7@�\R���.6�G$�:��i�m��Ʌ!O�jv6����!�w:5�W9+�����a��<T�hS"ڛ���]/�l�����o?1s�o��x�M1��M[GQ����޶r4�º���Fx�}��\F\sW�X�e>�δ.SP��,q���!�N��N�ØUp&����kse�H��@x�y�������]�-�$ND2��!���`��ERV~�2�J\X9XN�b��VRH����O����k����x~��5"|�p�b 
��|Aý��[�����\����Ɩ^f����\��Z?�v��9�.�/*q�U��_�(��I*�A��>�����/�]�N>���u�$N��$�J49���A;m���?yk3�\�0:*G�C�k�)��s��^����Оߤ��[�W�X~���p�7	�d*R��=�  ZL��0tO�5��)ܱ�~�U}j��45�Z_N0��Y�Z���tH/�=r9i�3��7;ܽ��}�p����@�KTm*u@5����+B��[? ����u�c{���N[�&C��zJ~e�{e���dh[k�Ѵ����fљ*��)��Z T�
R7ǥב7��'w��p3V�7x���]�a��k���SIPVU�o�g��a�L/}�o�?�Ka �R�-��`7��7M�4"Ԥ��?p$�%bX�?���T���jv�����!� �Q]�~�y���^Q����x����~(�;u�]R����T�d|,���������#ص�A�g��x��ǅ��R.o��ȳ�6ܝBoZ��T��s6�EDݲ�$����ir�l��	�R�L��]4��(��p�O��_^,��ND�X��2�\D�Y+VΝ
3�K�����8c�ߕ�M�o#���gA�%��xV�h�x��V���+
�|F�*DS ��X슥i(i���P��U#�q�a�护
��A>�M�A7ӊy�%d����^w�5�"Ƀ�/H�͑�<f�{ɶ�QJ�=F�i��������0�S�&��S|�;^[i�h�8%�oT����n@JA�T�����%n{��*C/l�a1���.�����@a�yg��zQ'�8ns}���N�$s�\$�xlC�5������:%�x�6�N�5��RT�(�p+`lK��wE�fU2W��G�S~��mF)?H.�Y,V	�*gXk��C�ͪmo+6���Xt��r�_���>=/K�Aˡds�rs؈��I�R'��mh�0���wS���o����^/"Y�j����ί��#V(�"U�\;�9{_i��#������Y�l3��|�)��Î��U��Ȭ�q�l�08�K4W���:����8�)�;��*���./!
�q�΀���wȀ��p"hi����jn�:�%���`>�,VΙ�ejAx,P�Uy�W1Y��^�	���^�L�7���PPo_b��W��Ur����HϦ���7g����Kʹ	�!���I�4�Č�3�.0�4�ְ��/apVv��{������q|8���z����t�:޾�E�a"+*�*�GHPx)݈G8̜���OY�L�Ȣ�T���2O�֏�ڏ��/Ú%l�*�D�E����ǀ�	L�ʨ�0&&��{]�5(���ʱ�PKV�������W>��h�:�:��l_R��j4������&[��n�/p]&%�x�/��1fwf��<']f�H_�����U�}�;>6ge�� 4�Z�<��z�#6�6�T*A��i�b���)��h]�ih#��}���񖩄=>�a�>b]乎^�O���8�|L�%]��mP�(<��aN_:��虔х3�u�c�T2�Hh��:mo�b�19�/>��[H���N���?#��[�½�%u�Yq��G�vj>i��Yr�a|?�A�;@�ˑ(e��|	�9���1jFׇD���&C��RK��"�C7����w���[0cQ�:Ë�ى|'"R����d�&7׍{tnްj͍d����X�U�:��̀Һu����#�,�R��������C�-��xDn��*�~�f<2���(����FC$��u����4�(i5c���\�B���G}�+�ͦ�l��yi���^������gB����X�{뽞:y6iЬ�5*j<d��5y��G��~ ~#v%���G=��˒fv�@AS�>U}��n	��Y�ҡ�+@���d��KǞ����G�gIrP�G��2z+��ʀW�거f'�J� ���#;�1�b���� �>���̫�������! ���T�ڴY	k)�K���)3�,��Ӟ��A�g�C���q��~ w��n�x��;�*�@��@i9�Mc4$�����+Fsӎ*W�	�7K쐎�n�a���vqs�>_o��ukN �@�#�0�E]��qд�t��7o�2�(��Y�?'��u�n� dx])����o#S�
��[�NT��(���ѕ�筠7;�ϳU�Ds^�o���FQ���T�kc��m]�g�ӎ�C:���MA �Od��n��xs��@����=W�x,H�@�A����3��C���Io �ewY0}B�"�bW#� UBq%�<%����/K(��ݖ���(�����:�|X�1>˰���u�o#����xq�a�UR.�b�9щ}A�8�� -��yv������e��y>�ިo9�ie�7!:��>��n�C��Ju�6��
i��(B�i�b���i�le!��Lq0�
-`�+�����%_s���O���%U�%���b��]c`���N�+���׶�J�xk+va(��Y=&0^~$�M�rgXm�O��bԗ���U�;�AG�j�9��Z�W�0�܂)��0g�٪]�l�W���R��K��Xd5�DV㳮,%IoeY��?_��q�n�|%\5���^�R�#��:�	p,3�>7A�Z��1{��5/Hd�ܔ���*l���e�,mw�!�ΟI�\A����9����D��2C���F��U�̃jp[��N���C\�����9����^�kt�����l0�ֆ��@+�> ;����s'N�4հ�4B�c��2���dvu��0fE�s �C��z37>�C�^��s��s�F�H�ͫ����M_�=�{�8��?`_Sdj��O\�6�Q���Y>�Nb��C�m0�3�
oF�w���4�TÁ5)��o#��{`�|�t�����ص��m�\5�s!�y�f����y�IL��H�-ݣz���N@�j�#��G�YY0��YحЀׇ����e�P����z2��?�nWjb����f�������>����d����N|�NX����WG�����&�OT�f���+�r��9ʙ~���~�uZ�!�:���*z�{�e�ً6�-�j/��n�i]1qqD�z�j��{񒿺[儴	7~Iv������������y�) �H*%��Oe�^���z�P��0�!�\��dD"��>�)������9ڌ�&TO��W��(�����Ē�^hc_�dxm;p3:��=R��m����v��*�񑽺����f	i`��W�(�_����.��@���'ou��z�~�����h�����Ű����Ir7�b�Z�c5y�MP��3���D.��,A��4����j��)1�g P�d�B�{2�s+�x���2!_?+zt��ds�2����p�r	T]������f YtC�tQ�=�����,�T5t�sSR5Z;ܫ�Z��I�[�G 'pK��;p��P��hd���R1�B5�m7�X�l~���I㩌#��y�tv�+/�!���s?�X���x%�@u���k��?��W͡�`h�JN��Aq8~H�u�q��q�զ���܂�����(X'���q�[@�?GS��^�rQ���,�TxK�b��雠�yLZ+@�P(�2PK�`g�^�(��=ٽ Q���.SnU��{�]��9��#��{y�,$���g�t�̬D� )&�Af�N��q��>�Js"[�a��yQ�`qK���	r0�h֛��4I�9�{\��A��E%bzA�	�+�ƽ��0���I�Ґ	�U�o9 �Dг�̬ߨ�5J�-��Kz<�	���:c���g�b(d�	���"����ZE�vf��+fڝ3}+�����}��	�b�3���a ��. M+W+g�j�n{���$��9�j����#� ==]���l��#�;vgz�	Qo��6݅�7���,ݜ��8O�nn�<]?n ��5rUoj�σS��#6��o\1������@��д�%N��Nz�>&S y�jTRU�V��� ��� �\iu����-^$qu�ST�l>7椧�:�;ط���&#�^H2��@��������H�i�L�;�E��\)�wЪ�.�wK�x𚠝bsc��l�$�`[MP0��mO�ܗ k>HI�智�#8?����.�k�~�A)N2�p�b��摖yp$����a�J D���1�v�b��m-��l��UȾ�d�#S�Cc���/�I�5c��p���ch�6�4����<�^�˙�uM��T�Z��/��л��62n�f�W&��D�X�x�l��).2^/� �B��Y���Z�<��ݺ
i-��Bh�;!���G|q���P�}����"9t7��<'�,X��l����]NܠLd(4Ax���K��(�t�V{�R�ӧ�����Z.&�?��� ���Z��CׯI��6Z��F�P�+�6�����2�T�� 2�4��~�(s{Y���B��Z�o�J��JL��o��\k�%�3�7��C��1��,�lZ�u�����L��w��_NH���ǽ��nC��!�ԅ!��f�ֲX���Z����j�e��2���3E�2�{改6Ya���NO��Ć���i�=����}�u$,z�"v;${>a�|��j[Xɯ?��.j���M}�*��j�E��ڒG����٫A*ԨЀ�Q���i�y��`7���?���E��I�d�u�� r���	ɫlNF��t{�z����M�&3�u`u|�ߚ�Vq�-�$�fup�I3��z3-��wN�@<���I���d���Z!�;U��J��%/r��6.��7�����-�[��l��=d�:��_MA��V V���N�>T�3@���"�f��Yz>޶����r�+8�$gh�Ў�3)� �iD7�"�dt'��.:n��$��z��nK��m�V��
;�MN��U�![��8|w��qPr՜�2Ϊ�v�Ϛ�_���ӭP���P��6��@'B�J��5{*�챎�R��)���-Fm��!������OǉV�3b+�xS%�Lt��(�$``V�� ��-��A���Q�?�v��yL	�ܛI~ �=s��n�3Ҷ}�ac��s/_��O.��c\kP���F^�+z�hu}�\:�>�+|=KoCgDql�rb��)W3:;G�@�{��g�3�[a�Z�m�s���VA'�����{v�[���C��Vo���L�����5�n�i����c���v�aG�MC߉�:f��;�{�]�&�7��uRiu�P�;[��3�#�Dy��ȉWI�KSCW�����R���+���.Мgy[���; ��oI���A׳b��.]�ĺ���$L(��R0��� P����]4�k�bXa��=��#?�m�¿'��;*�> �t|3�\�V��!m��Z��fr[����^vܗ��v����ً�&�%R��'p_�����'jˊ����AO�s�ϫ��+�����@���2cKl"�/l���-���[@UY�㒯9{r�H<�g_��nD�uy��ț���ƞP�VC�2
�}c��`xf8�]a�B\�F�K����-jr������u�Z�#(��Q�d>[Y��M�%�
c���V��+d曈�i�4!�n���q-��C+ff:r�sfmuX���A��:��;�9oE%�+�Iel��@}�UW�ʈ�>��W��ֱ�3ӇX5�\�ɴ͡`e{��ZL@��ن�VӼT(�|G+~|�p�U�Q�wlI��ح����s_D�0�����/$�G~ͦF0�RB�\\6�=yN�����(g�Y��R����V��a߲}�IMG�&I����L<�%hlp��n��uYS��U�]�'ܻݹXk�(��x�)���R�����h5���Q[8��P�Y�J��I�=�jd'9�BP�t�I�ڂ���>��"	9� ���$W��*Т�7.jms8����fw����>�y!�Y�๏���U4���F���.��>"�����y��K�����l��� �9�ԍN/�Kq[&du�����o�0�{��AU؋7�=�~-����m:�g�	�*L���v�������W�/�|o. ���8��������?��
a���Z�ݎN�aO�U�Ú�F��R���A����I���{d�w�J�N���Ŀ>,E�����pʑƩaѥ�ZY�{2F�%lJz�s����uL�@4A���	�UA(�-�,|��jL��i�~o��	Tph]�32Y<���B�B8-,����f��\#��oE�y�+S"70� 9����$�]n�?�9��_�� ���x���^Vyu���7��g��)5�8^���l��mn'��|9ݥ˒�Q��2Rg��}j�����H�	�њV]1���㍑�i�
�d4���{�*!X��ڎ�bW���!�݅+|����*�z�A�EP�@A�)J
MM�Z���#���r/X��.^���(:�A�+�S7�,���*R��-����P�@�d\/یJ=���l�qP��\�꾶�ɤ��7�^�8�u��9�ו�Y���r���ᦣ��Py�L�b��Y~қ�#�f�� ���,�����6)٬�:=�w/�:���;�*��OOӫ%r��1�|��ڃ:Ck�瓔����y~�'��'����Jg��`��}�ݪ2�op��&�t[q�8�zɴڹ&���۰E��2�}&�<�n+1��,�^����M�.	�.�?W�%fډ!u�f���yjO:��%�5��1��J>�y�^�fN;�+-���/�0@��m�-� b`gW��-yW�!�d�a����<B�{e�R��V�V;�[ Iă�2�����+px¦J��o��I�t�B��;6M�F������Q�T�fk��=�������&{�� 00bk)����n牖�B����wr���2I����9��\��������q"є��5K�h\l����v�c"�C�o{p�����x�e�����m���Zz<�;e{9E��r}i֝��}�qj@b�âI�2h��ֳ���{�K�u��G��άyP8����L��2��(GsAL8<6cjC����GA��RX<2����H禃g�
w�z�MYf�s�)\k�S<��R`�y,q��aғ��c]�&���u�+����l=�o�T1�9m�hT�IDk��3�3���{�\e~��fY���{��,�ɛ8�י�(�a�� ��?��_��;�z��0|ء��V�����vgX� �����`��+�E$��?}�� )o#]���M6*W��5&Si��jr�|�B�by-�w� �6˿w�����~وy;�v�V����m�'�0oӰq�7$'H4��T��O*[Ǳ@P�F��/��O(��zN\�⒦B�X�b 3b_ Fx�.^w�lWz�k�� @[�V�P8�P��[��M��`���إi�]2�{����~!�i���}H���N��`wm�L����)�!�)�������ua��7kZ�K��]��q7�|��w�KfPm!}��Ԕ�jX���%z�Y��`��<��KO����F� ��~�-:�i�I����ns��R�
�\Sú���۹�"3J����mf>�j)�3F�(��=���\�>h�j��a�_�� pH�Hw���0
���������t���:,�7/���+ʶy!��Sx"Q~��6u�V5쯮nQ�LΕ��zI+�?�ĄQ�R "R+��"�pj�?nh�eF��������6�������,�
��oky�ï��k�A��QH{2�Ƹ�����-�$��H�<?��L���H�5�d�B6T��UZHXG
�.�З�i�Z�͘٭g+�J��O�`k˟F>�OS|�,5#����v.���y�j�5B���T��XL�w�7V|Ǖ1�-��Ii�l�9F9�b �H�w���w����C�K��ك,��yc�7� #u	�`  }F/R��p]31�� ���rK�<�g9��ƉQ�H��OՖ�-y�ۓ����_	�s�A`%᧣ph�;ב�	�e죫��vz0O
E�����ZA��>���>��	���4ྡྷjf�`@$�>�ſW��ج�.�� ��JZ3*��hj`�`�b�2F��̘�80�W@�݌�A��1�'¾w�R����X
�vD��ՕkA39.��#h"�f�_�����W��`y˦v���k���P]5)~g5As�����T��K|Ay�:1$;��Y� F�[���|�ˁ�*��\ҊH�f���n;��wU3+A��s����Ѻ`ȕ����,�e�YȤ�K�͕b�T՛ *g�ę�k*���(va�%R�Q!D��K��0��kf��Hg�K��>X�٣��u�u�ޠ��1 �2p��Ϥ�*���jҼ�+��Y�42y��0[WQ.S'J�%�#l#�[N胄�D�����7+�YC.7a �BO{�ȣNh�]��_p�_���6Z��¬�IDᜊ*��j+�`3Wp=�x�R|
6�����B~!�������Zf�!�).*vg���ǯ� �$���c�!;V@9����aA��cɘ.?�N���+�����*���Shۗ���~����V�5"�ꦓ�me�Q�գ,�T�s��3F����(��3�"h��������H�E&i��	�����BıdqЙf���G�=�V�y�#�`�#�Jr�[�v׷B��*村�=�s�4��w[�=~�eS��\���`Q��k������rO���T ��S�3�J�=�X��w��jz��!�6�?��¥O�P~��K:Ǻ��7�A�zJ$��~g9ٓ�}Y�, �(x;��t�pD���w%.L���]���j��b|�T�U��#�]�q$�^"�����~�51�Ccd�W�v��#�Eu�uD֛�6�'���&�@�t]mH�i�zt�jm%�:�b�|���!ͬϠ��~H�~��y�P���`�o��1ku�ɰ��`V��W#�D���Q�ja����W)F�V�AG��3�ղD$�ҸL�pE�qJ��>&2���t�Vt�s�m��@���4R�ח�4ۻ����?P��6��CR��W�/�Ǣ+b�xRnJV�L@���pkK���D��7L� y^P#�ss�N��Q�%_�N>i��I!�v?�o]m�Z��E��\w̌���!�$�{�BJc?��xb�~�T|;��q�1!=�Y�~-4������KE�������{B����PBv��/+T<;mCgU����Rn��̾c���ooEgGC˼���,�,��u��H�x�w}��^zͫbѮ�c�CY�(����.���o���~��07�!�$7�ۚ��غ^=h�LE�;[W�.����q�z�Z�h�2 ��\:o�+ԉ�F29��M�d߃�Wu<I1Ij�Q?���s6�{�߿7��.t0��2պE�%��"3��a�Z<���b�p���d=Hd9Ů�y->��^���6��Ӱ�cK�O��`1����et/�����bR�'������3����6�_��Q��󦍬�c[E?	h���;a��w;�E��&��F�T�m @���CHO*7�ڍ���c4\ω�z��j[lI�@K�ƃu��p���V["Ӆ��59>��a��]����3mb<1;cߵ�o)�cވ�X��p�#UN 4��/� w\�`wLX��h�D�xb �_c�clSܠ���L74xF���a�&��-��93���a|(�f�,���r3�s\}�!���A���=D6\�s��1��,�k�i���4ޱ�W�?&q�l&�T�x����Q�LGW"m �)[�,n��o�M�H�kV��uk*��&j�����5 �����+�=�ַ��Bj��PmΙ�+�A�:b�	uX.���ڋ�y�	|�� �̲������XY�5�5i��p�8�a:��e&���u�c����_$�Nlf��M�հ�9�A��c��ZDD4Qy���\^�ж²$���U�U����W)~[�^W�[ԲҲ�s���N�������'�`�����
�k��ki>��~4{���?Y�W�:��`$[�b�#���1���wwU!͋�[B)����)E�o���ߢC��I�����mKP���������W�j�F,�G&J�K�Kc7�r�Y�N�t ��ф�#kv�#�k�j@�lV�+�>�x�`��\��n���"\��@��1(|�������%7��~Ո��%��4�ﶈ����d�����0���I��+Yu��J0VP��+�fV���-��i�94��,�$�\\BV��r{r�J=w��[��y�G$��_"�^�̞�,��b熚m�U�=X�
;�x���BUN�������Đ��ă�����(��Ǳ���#�0�x��B_�C�D�6ʞf�֭��Q��Gd�	y���7��W��1o5�����	���{42��:�1�����8���Hޓ �:G׃6�\]�t����boo��-��<�����*�����8Gc���%X2Q٭����- ���
J`2���`��nQj����^�!]��/�	h���M���`��7�}��MWJp�ɒI�ClLҒ8�Eʛ���0�7Ο�R�k�/�4��y�R��Y�^�>���_� ��bUk"E��~3����H+��^�O�d�0��w�8���u�����F�oU�ɵ
WW���a��ͯ��]�6f� �*ث�܌�P�H@� 5n�]eg�o)o�7k���� t��%Ť+]P�䑝�hI%-�(�(�HDRP��ot?8ǥ}�5�l��fN0���,.%@�r[��ǌɔ?R�Gk?�W�gF����-��"#�
�ex%����O�B�쨠���&�+��ܶ�����5Cq�X�W,X�qX3M�����X�7eaɴ��Y,��k���k�ϡ���8\͐�W�E���F�i�	��C�4�,�e�`��UB(��s��Ã �*�d?R������������$F[Q%h"���Om���AG�:��N�	@U�6�r٥���[����hƞ��>��ϺP�| �W��;�G��"�����̆5��s�ʹ���taY+�gh�d�鏿��`q�U��]��(�?ACAU��]B�>$���������ς&������1OI��uY]�3R�մ*��A5��7|���m�Y�4ԋf�4��}ߣh�[�W�}��g)��B�:7R��<Sd�@�N�o׬�H�0�qv��r��]�r�(�8*��SH27�8��n<��ɬY�ӴdYb�@���tӽ<���Ԣ]6��YX�1@�B(+H.bPS�R"��Ң��{�]�)��o�0���΃p�K�a{�z�x�+� 3G���V�˴N�?�@%�;�qL�a�E�pj��Og{��i۞�<Ѩ�K�8�s ��>W�?�}�RL��[�o���1Y��LZ�� ��ͪE���	J�����	hFI_M�q�g�Z�Y�m�Jn�+�{�4&k3I�,��P��5vk��B�N���8e��T�,PCa��P���RU��φ���Sq/� ��������[e���\�#9±��`��f�\`'&#���1T\��"�Q�ٜ���& ���9��}�ܫ2�m��O���;Ȏ�Vl��ْ(M� ���	8s�j��d8���bW����)jU �5{{�X>4�9���>W��z��saU��|�}
y�9pypѻ�Tdh+����*1iVGT��ܪ���z�~0�2����Y��s�S�]�' �q� a]�����0v���Y���]�N|Y��@���T�;�J���o�E���=�|#�퀳݆��U�6t ��'�S��4�$��#�#���}�x�/teW~����e�#pq���5���V\�O��[����v���m��A���r�Ӧ̠Z�c��&�ɰ�j5YX|�lu�5_S��s)ο�N&Ga���0�!k�Ñ:���89<>mL
ALr�+*|����Y����廜������LV�^$�O��ow, #������c��L>���-�I4&�����&Wb޶?h���6tNB��
+'6�Εc |����B�|�8U2V�� ._��b�c��q�<��%jȮ��6QC�2l5\�I�zk�=RC���^æ��J`)f��Wf9T}JQ���j��B*{cA:��=Ƴ�jH�RV���!:��&ܭ����� ]�����γ���e	�ٮ�(��2;�m�I���)`�ѥ_h�ɍVt��E�
�^�9䯝�	F	ZF���ˌ"`sz��D��� ���Nd%�Ә�˗(>���[�b��]�z����"�=@NV�J�jn��&�xL-�(kMe2�|g�=`2}(�hq��bx�T�3��7�dP��٣5�aH2��7X�BX������6���O���/c�gI'X�&�w��S�}�c���?���*��?�SU�pq($��_�O�Q��n�p'Zj�m;��Z3vP��� �ˉ��KUrP*���%�]l�c!F���hMV5�c?��TEo���`�"S���E����qa:��Q
{Lo�$��cb @r�ok����׎�2���y)9?�N[_|���dS��w�g�>&����m q��Z�Hؒv��0	դs�V�k� ��+�Y�=�W�u����ڂj��?F@��9)��9��<�f��a���I�be�1����&�� �u�PR�xv��/������|�lӹ�$w��� ��ld�,H���S��[k_�F���_��p!Y�!缃��!�˃��E��I>��տ��V��^��mp��E�+$5!l}�z�x����}1��=oK �\����e:�B�E��UR�IS�:�����M"L38�0'�t�ޭw�U�ݹ(���L�J�C �M��e%���b	��[��ڝ�˫�%�e����Ҩ>���3uӏ��?���v�+�%�PX��J�s�p�Ob�&C)+舽�mAL�jϷ>�b�,Z)H(��״}�ԭ[��|�k.�jpѯ#�B�;Kl/�8��~o\���-9��_8�ɧbK�44������7��$5��3�O��@�����;�)�e.���=J�����S;��rW�����|������D� =,�G���m��OU0/��R.=��U�{o5�ݖQ���J�%�Ԫ��e���c�a���ͿH���X��8���hl0P�'���2�1�����p�����$�XV�Z�Jo�3����Xx@K�r��汲8���F�ˈ��/�,��؛�:�~���9�Z$QP
R4���_��x��`@=�3�T���:2~�%��	���c����ڼ�/����|e表td���(�p}�	��aƂ������L��qF��b��רC�j��^G]c��Ҋ�c����+�]�����L�/)�($:�$�"+���R5�g��Kz&�Ѥ��=� �hZ������h_	�{B����)M��^���R.	@�qyċ��UU��[�����q��Be��V�`;H�_ �X�\"�2�: �$���en�X�����#(Y��Kt�/f����K�T!��0?��V'��wcÛ���^|�w�8��<R�<�P�p���O��v����ĔHz�-~�$'�kG�{�Ҵ�Ɣؾ��V�<�Rf�$�o)7&��"c��Q��H!�m2����O#BX3R��Дވ�σ.�_oBK�Tdo�4�uJ�]��1fh�{�$��C��i8,`��,�������āM���b��������O���(m�7����Z�ɒ�Ra}
M�|�h�g�b���m1�I��x5�&��{����RTy�B=�s�t��T���:wȿ\�(����#��Um��I��iU�Ʀ@<!q��
X�)6���UMqkR[}&Zr�*����W��a2������P#Y����،�8�����&p�h��B�ځ�u���T��?�`�����k-���A�}�ׁ�B��w��7�I�w>+���U�6�4vC�Y^ц�������N�G6cJD���(\�<�kR����]�b���e��<�"ib`?���m����SI�J;�z��U��O�cdPs���^	��#^mn�*ᚑr;���WEꜧE��R��?�=�ri�Fq��u,�$�C�]����H�&�6�������~B�+� �Iot!*�6��ѐI�g������2�fT�m�3����&WS����y�V�����׸z�	=��9����o��"��9ck8I*�|i��ɲ�\�n�ԧ�lC����(pD����N_�'	j��r��~V�C�C�Ȕqj��q�9i�h����X��~J�o�ZAQ+g�9����h(��\������<�M`���  s�D+ �]7�DL��C\��o{�Eb9.��7����H�.�h�?���)�8�9�7�����d���[��F)�%�=�F�+�H�Y�˝��=_�� >W���'&����c=3e D[$����(�}�|���;A�,]m����T��A
�(�G������;��;r�)�l���b��$���P=�a�Lh��ƗUK���e#�7ж��"�O4c���Hb>��~A��o&�Fp�����Osb��V�ϰ��w�Ie�I����3p���z�3����:�h,w�r��'�K<���s�&�ͫ�nlY������В�bn aU?�M�R�S���.z����M��K�J��D�~�EN�ٟ*��=���L�ֱI
y">�O��x�����s�Qc��2 FӮ#Iˤ���~j�-�Щ��N�w�r�=/�ߖ}�vo9\�1\��v�cgFCcS���� �^�A��a�������f&���H��>����pȈ�@�.FIu��]׶�%6�E�S�;B�ʴV4��%�{6������<�U�o^+<K`�/ʸǩ>�2,?�݂�=-ܫ׸��,{��Υ%uQ謢DQs�����Y9O�妞�W�[�lՌT���"��ِ�e-�	��`���GXni�מ�����;������'�񙗠���Y���\P�>1�E0���'�����,��m8	ԋ7�L{?�����2	@w�ĩ�4��B����<JpYx�T_�!���^2{�[��GBD��x+ox��"H���#����N	��3�NP�� HJQv��V��-���Â��%���M�wD���A��tt��=�<��ry���ͳa�#�Gp%1���Xўm�-�h��D�1u�M)��s����<k1� UckyO^�xS��ّNSwC�"](G������O ���;$��j� x�_2�e������ޤ5���}�,�����4N�/<1௠C+\W3�S��eFIa���u��y&�ŏx_���DeS%���U������n�3�@U:�@������C=�l��`SϠ����c�5�L�N⛖"�vg��|;G�d�28&t-���������,���s�d�j�Λ�[/�&�7�,*����Bn��I�x�B�������
��փ��$,g�<\��4�~~`�'��F�9�\>��M��|���Ԝ�_��k\D��Efŝ�u+R��&$-��uv]Nz�/Z���+٦��Æ홰�����p�u��[� #�(.Y@�a
���9H�Ek��q`~=�Q������?�߈����ڡ��3Ѿݑ��u;�[��懪��z��I����U����&;��K� Ao�e )Q��H�/V�뷣h9fU�O���=�>"N_>m�����p ����Z�]���Ϟ�m_�NCg�b������cl�'�������;�����)Q�D@��zx��=LPU���P���6��n� ��Q��u>����>]�^��g�-�e��R�1DK�Jh&�,�)?�8���L�4��llYʹ�h��[��mS�m��#��I����e��l�#�ˇ�f��P����q�1+/�����͐г�g)]{���z�!m��p�\�+3~2���0����pmvS�v�C�L�o���הs�)R��̰��im����#�ALIva��ƛ�����3�=#.b�o�{*@�#Y�i�x?(Ra�����t����x�ql����t��$��-o�dM�"^4l�լ��T�M��d�eQ5�~����M�v�ʸ�VT�h~qrD;��,F���0hB��Q�E-� RD�\U�4�k��%���۵�o�����g���� �NN���J����ݼ��zN�qy���B�1th�i6��L<�ϟ�鹣f��K}�=Ԕ-A�00_�?�!�����Nn�0�>hU��E������l���� {���e�7Ҷ���g#bt6��P{�`ܵ���,�/}�����2� 	�w�IP;��gr�U�Mb��V�GC�WE��� ��z=`���%g�h�~}�B�H�� ��Dl���R�%��Y9~�+�ѻ��`�7��W��[�|��څGȧY� :��.��eC1�O/kA���K���-Fx��E#�c�\�^d��%���s���*����{5#l=�=hfw�v.4�u=M8+����[S�)����W�!��Д��D̒�3<�2�`7�4��zy���QMR��uM�[a�?F�O2��-���A	\v��⶷y��~{��9>
Bh����#����
u�,�����a�����7	+'��k�!���k�V��ҤY��dNv�s2��QS�+�qk1^����Z��
9�%cJ��}p����-��
\�HP��٠N�냦������K ,h�剘���q�c�}��_Y��2��/���z^??��{�{\Y��&�TI���S�3�^���b��8� z!Ou������0��g��㷂�j��������Qָ~i�jP�vWT2W�þ�=�_Q3�":�c*Z32.�.�vp�fq��� ��h��vg�r?^�n�q\�3��~����%��AadR8,�gΑC�
�=��w����%�K�P�����|#ӉLU!x�m{��|,pu���~�Jz�����ATthO6�o�-��
XMvp]}Ygκ�
�{)ֲx��0.j��4٣�v�Z1���q��q[%���^,$\ϊ���n�p	�l%k�x>ѵ�[m���#��]9��#?+��GzǏ�����Y�^�[��q"t���̯&x�y�@�6�FhlsW�|{&�}I9A/f4�5��3n��)���~Sq��������W��u�q�P�.h�]GakS�Fڡ�j��w@�g�\P���I��x��T&��,^�4�b�d<�BS���_�D��E.č�Ŕ&!�������%0<z`��{�`��Zw�Y��iH��ב����/4K�Ѵ�G�bH�j�>u����Q����_`��
��SO�ā����=C�k��2��;p���=8Ѡ���=��(��$�Ӟ�@���,��`0a1v��lg_O�sN��%��Y��~q\�wF.`:m�ێ�xd�ZcB�_�ݢ���j�es%���q��5�DNۿB+;V�E,D��Ě��u��;�����@M=Ԕ=�U�U�����F�~�=z���5:���Mv[��NmѸ��A�c��b:VQJ�Q�} *f��d4~i����e�Qсjb�cW�3i��aS�-��j�䉠�Ǝ��H*C{ąfބI*����:�֐["U�&��f|���MV=����F>��n|6��#R�'��ʱj�D�y)��7[?ن'�l:��F�Y������9����N�<�4]��]�_w��~Z u����㩆�P \��j@�TV
�., �?÷���s�=s��\+[��2��0���4Έa����nt*c�7^�!�q�/��j���(i�U$��M���`і�>x�W��f4������%��n�Ě�[Φ>a`6�$�k�;�Ρ�|e}��sđ3�#��$J�lO���� �S����������BBt���֥x�|�<���(��G��_V0Dc����r���\5h�XƏ�1�>��Wf��yQ����}]VI��K�Y�!�$��aW�6���82���ϑ�6" �nU�$���\7~"R�ј���P�`۝�>E�!m�g��h~N�0p�f�*b��*��_�h��C�TW�Je��u�+v&Bܒ-f}A��鍻���L�F�M�L9$��?qy�RC������X�����5����}l��-Y�s��������տ��9p�|`������������!�<�,\���1"Mt�����0�'�*p4QD��`�ƥ��\ۛ��v��]��>��+�]� sXX����a��M��6d�:��u����p��:*)�|�3���k�b�I]\�,LSG���� ���5�f{�����:���Bk���kG�5�����-�{��m�����v��D!Y�-�i@iBq}����Ӷ���ѧ3ȡ��`�zY�P�G~T����;�O}�m0��Q6�.���ژ	9v���)7*��U���z؅��i,(%e����d�7/}��c��S{��jأ� ����Nk �0-x�bН�����B�o�����v�[�}ٖڐE�teg�\�����4��$=�~�ªÔ���EK9�Y�T��܄CjqИ�נ&�0a���ǈ��	�3y�횆��2Վ�vɴ��9@��;4�@;�έm#�m%뭔��N�d�Ɏʂ��f$�[r�6tx�����/2�Jl�ʴr̔�|��?�[�Z����D�G\�$^�����R�w�h�W�p�5*s�ȧR$[�$!�x�N�\pպ;["�H��큿���nk�{�1��� ً*�W�����A��Y�c�kM�]��|������d]o&��%~���D?j���F��G|y��N.�� Y�M�c��8�2�rf~E�C�M���n7O��cNH^�1�C��[���ܪgL�3ľv�Cn�s�i)1���`]���*��ה��J�TYcd_���ePP�Ι%����OHqN5�#!��X�2�3SCm�J�~p2K]�3���/��m�i[�
H��c欶$�e�t}ICK˷!Ϯ�$Oj�q�EM��6F�<����/��=�F�BU���VA� *����92��dMjmh�f՚�t��: ��>��"��0�͒{UFC���>�tw�2�oI#�.�_�it�ot.�D8Ok���+;�j�	���d}T�p�E�;�~4��H�Vo�d�ƎX�^��V3������*U�����B���A+ ��6'"�{�|q�̟l�&V�+�v+��!YYft�I��=Q	�-C��K��r�p���"��t��Sar��E�zDeC�Gu�c0��`C.������>����,����	#	���dƥRr\�� �G���=f�?����ES�F:k zE�`[�Y��e�$	k��>���6q�Au�_��차��vJUAת�����G����.��Lc���l槺��k�27.A������t�S���W��e4�]��P˂1 ��b��|�P(����4Z�+&pIӠ�����S���x"�*4�?��8���Ν>as\�d�\�q9ʏ /ܴLQ����T�C� �G6 �;,�6T)	���;��j�-@zi-���c�X���<�Q�z� W؛�@T����b��>Pp���}��5/f���|�z*����F�F��\�?4;�gA��o�af�,��{[)�~6u��g�O(ln�\�=&�I��^�ń�w�s<����`*M�K�T��� �*'|���O���5��\ �\�^o q��)���]���W@�A�S�^��[�l�F��t�X��<D?� g�3���K�5Z;�M�It�Pw�l��
L�B�R�G���v묧�.>�"���L����f���i���D�տ?d ��W��VY�\s����;�n�,0�����a�AE!L���3x	��v/Q3Z�f�J�]�HbQ������ ���$�vd\�k�y�7@c�"ߊ�������1��Z��(�C�|�db�9+�����Mj�����n�KI�Mg܃�D�I��Iƴ	_�U3p M�'���k�2��N嗉U���~�\xO4���p�5i��;;)OU�5G������$G���6���H}	���H���,��T�mmc��X� '���>�Ph���Ҏ.N+��� %�uw	��-�M��T�:�}�0��B�Ȓ9595�CԀ�M���E��>K��kytn�hr6�)��e����R�2)��
��c?�+oCt�C�� �ڕT���4p�$�7�9�d�q��rBY֑���e��.�Q�D����ֶA�,�k'���vgC�xa��J&Q�>��lm�C>�NS��(⼸B��l�0s�/Rk�^�@^
,P���w�%ی����z%d�-���D�=�a�.'d���F�h����b
nxG�$��(Ԃ��NzZ%��͕�U^�I��#U{du�ӧ�[*_Q*��8�oIې���l��8�;�:m����J�&�E��XC�	��z)��jb�)֕�PC��O$W�x�L|U�o��5����,ҩ�4af����h�(�,PaD��<پ*�ҟ����̱��*��Q�N!�"��?�N#�
Q�����V�8B�\_�ʗ�[g^ ���u��\��H��Χ�g��N���>7b�����j����ӽ��9x4�:�L�[-C�=�\��Bg�U��#�o�
�S�W�2���E�\� 8d6�.��`>�R.�"��{��K��//S��A ���_|8qȔ��2r�s�#�����>�s)P	E0�)+z�QM��"F��5]y�Yg߃P��+�m��`C� ���>vh�72��"a�_�������c���P�ɮ98��Q�g-�ɣoR��C�uͥ;xr�44W�m἟����s����9����uXRFn�ڱP8���+�`����xͺ  �B��9�P7��`��#�̼�2��i�Ѭ���)ĕDB墌p'�:��Kw�`(�"�Z:�_���Wݭ5_j� ���'�R���s׷�9��cZ��+�Ͼ>��*ë�4���:	���#Ծ���(�!����<y&�/����W[r��>��=�:�ʑY(a��D�c#ۺ�t`��S�R~��,�de�3/LH}�U��Ԍ��i���۳ҧtn'��Gy}� ����:�ZBW|�H*��8�$u�{����h�'O��˲N��|w�|"�u�DH�P�����̫�[�?�=+ak�I���շPR,�y�d�_���Ҕ�U�.��3�zy���&��TA�,��T����ɍܰ0"�V����c',dx�%%H!+���Z�-隃ߜ�C
���r[��
ü.���J�[Y0)#)Q#��5���v" ��~�)*��a_�U��Dȫfy�TS��wS�x��>5�I�R��U��k�)���$��AYu�r�����P+%ٍ���#����f��>�Ҷf��r k�(���t1"#�`�SAA��4��� �������S�h-�e��MSɗ�M��pUتtV��t�2P�逼ǋ[Li3�c�5���%�����\��jK�e}a���V|��I��e��E�~����sC�J%����� �&�5�P:=c��()!F��M���O��;���Q���Z�KOt.�6HN}1lp��Q�!2��^�應�2�pg�й����;$ ��2wœ�"����M�
�c4��R"��C�BϏ����P��$�U���1�w�dPR:�ɞ��I���J+?���z�E���ӟ����\��t�J��J��v�>)�֒�C�qcs��'"��pa�9�x���;��oQ����I��Y���Ӣ\(��f�fI�m�8���G�՞����N�1��/i����;�Iw5�/�A��	{�~A}�9��{q�lۖrգ�����uR
��a<p���Tת��M�ϫ��厃@�>�5Z�8N��Z�n7W�.)Z�e�Z��|�RT9��W8��0�_�%uPq�JB�K8!�N;B
��+�н��D���х��X��I��b�wU�������ܱ�x��U<��.�V�F ��Is���-J�W��] �/��E�3�1HA�WQ	�9����Z3�3�@��N�m�]���Q�!<�v����Ģ��2��ȵ�ȣ�S��1A&���Kk�U�H�c|����1���B�F �p$��tJ�Q,�1�%�B<�M�t rQ�>��j%�������.'��5K�#�ŤU-��2*;��IlGܪ�!91�)�dM�I�8p$s.asx
�o�7{A����+��h�V7��)\X�g�[*-`�ߝ����i����L!Y�ɷ��cEK�M��n������d�0�.\�n�P����~<�7?p�%��JIhG�>����v��-65m�6*@\U*1R��>�%z:�köPЪv��]�	��2����ims?ɽ5��<��o�V�K���G=.�R%����W���m�:�`�)ǜ?��~t��"�-%y$��	���]��Z6GzM�����y�~�z�wI�zǯ�ܕ��w��S�O��Pr����@��U�=��tR�r%�e���_�J}��r����|�s��K���u\�o�\�[���.�E��A? NG�Os��%��R۳�^>	wD!D���A�Xk���R"����\��<£��?�����!�<�1����]n7!䬖�5�enr%YuU�Y�zm�
�@����(�ZL�1�Ƭ�|]2w�B�L8�V�z/���U^p^��)��쐴(�Mc8�L���r�W�o�b�=�mt�ǣ3�KB<DSi++O�i1:�����%`��tƸSp-j`�����~ �5SqW=�}n�u#�r?�a��N�r��%�Hx5c3��v��ޡ&�����|���ح��_��J(����R���A�i<[�?�#pSqɉ�2^�[Pn�<�NFհ�K�'T����H�rk.�C�)��E�G/�F�r�0��)(�-&Fࢽ�`6�gE*j��(�J�
`����6dx��9^X��)anN�X{���� I�z��g�7��M 7o�'%�L�wV�5��NU_J�p��;��2��.�^F}���/�S}��+q���Wn$zF@�L!Pbѧ!=9A�m���ZJ�����ɪ%x�����Rʫݍ桵�w�R�<����4m�Ң��_�K��<�5�j����$k���s*L�N�M���� �(|o�*ʔ�&)���z�@���~�7�7�-
	x�ͣ0
sT�5�e�ZQݐ��b��	�C�c��C���>Rװ�h��>>�-�¤F�)�R�Tpǩ�!��XM�t���K�Vv6�?��ĺ��:b��� ������2�U?���)�t��x��3�f?ĨZ�}��J��
x�!�_m$:��S�#F;�~�a��j�Q�1;�d�8�Q��	9%�~�1�q�ou9C#��b�`X�l���yr��KH�ʌŖu:�T��~�����M@�&?X5UY�#�d:����#wI:�f�ht�$������|w-==�~�N@ƮR\2Gc��>�6�vK���W��+�P�q����A�A�؜�� �i���QjD�U��u���Q�r15D5��8�V�<�%)m[C��}J)��1BYn���mI�X�}v�dk$Ak�wМTѭ�j	�OO�kߘ�������Z�U��tH��I�?��]
ҍ�$�7I�w�;��PK+���d��97MpD��]g�CI-e�s��F�`�C"*{�E�eg/�(��4��o/�^d����L����X�/�:�W���a��^I��h1t�<�X{���9�	�c4�ފ�ǈ�2��ȜD�:Z���B7F����I���8�+Bg�L9<,qo皤��u�"��O���*��$��OP����+�)�v�X�*S[ɘ�&�	��/��&9)��Wl,�vF�[2�u*#��3}�*�Y�Mw�3��0q������j��$�{g0�'r&�J��*��9��#0��hV�"�9�' ��I�G�0g���êJ|9�%��ӳ��k��R�Y��O��\�?�i|b�z>��-V\2�i��)�n�2�$�2h;����s���`�>$S6d��0"�7�c�4>��}��b�[�Nd�k]��"��:��`�$����/1�[�m-�q��O2R�HeZi����|$�I�(�5���{�alP�>����8H�ف�yT�h�)p=�϶=�L~�U�4m ǩ����{�Z/RY8ߢ��k�%�̎��H�_�B~p�ܧ�%^T�0@dU��N33)�� ��u9A�kC\u���Y�2�Y�D��){ר�J�1���O������Ո�i�9���۞<�M,�h��?�ŘYBV���8���<��z�q$��|Q$�ޱg�"����+a�ŭ�`lr"�EI;��'�-b"@h�HHj�rM�BD��,�Hā�Θ�
X�KUҋ���B�U�=QE�ҿe>��һ�#�%�������o���.<eJmsm$^M�Ĳ��	���$�{�E�Z���~�p{�u���en�[����$�(䊧weӉF!��}��Wb���:��Q�Ahل�x��ui����gG��GX1���HZ�!ʒ�^NE�+89�9�"�/f᱙٣����Wp$p�����ܳ�pD��3#��[�]��Ŧcd�#a[��9(���Y�8y�E,�8�0��h匮,�-��B��%��W�7X"{�r]�W�A*@q^d���e<ْ�5{��3N�'�fg���d���׵}�)�;���,���d��Vw栴��_lh��N~TH�n�8���bu�PTDϩW�������A$�E�&�x�+��bg��'��K*6�.���^ٴ��Mr��slt,r�V�1�6���?�m�{���/�Ch>�#3�[v�ߵ� �h��d�:�Oñ(�bU����/�A��0p�E����'�%%�����Ǐ{��'AWV���3п�"5O����vKN�����)s�R�g�6Fׇwͤz!�6��oV�Ot"%�EK��4Ԅ��X`[�E4����L�ϩ� ��#�����~�u}Ϋ�fWI���d��k�e�;����F,����xv��ꭕ�*���d�.�'˫
�����jg	,}=����7�{�Zޙ/b�z��*;��d,&���6r� ބ�s� tix#���Cn*�����(�pr���&���wQ���x)����e�9��FI�+����g��!��u�+��Q�ī1!�׿ ѷ�T��k
^�N���#��9_��z)1%ڇ>ZP%��?���^-��f��3�~��ۺ�Z�{�Q��1�.3��PK�R@6G�N�D��wŸ���v��i4�i�r6����f��4�������G��9
��S�:'HLƫA�bx�;��P�u�>^�Y�:|��9�b"O(r�d㢦PƋF�Y�bzv.I����5V��e'�	�I3M�%���H�%1)Gku��'�c]f�6�ȗ����(�r��l�]t�Z�|[����q��=eͬ7�QD��Bk��
w�9�s���.�O�pK�85v�g�f7���è�|�0\Y�m�A��B���3��PT�D����r.�D��ZrBL�
m�#kWG���5���'+е��`�Ym�J������f�b�� ��a'8�ny s�D.� +ӭ]�3�0= ��T�L�*��l�딲�H�:��or�7p���W[�6����&k�	�l�}?<���ى,ӡ�^�$BA��7_-����L����W}"u��0����Фߛ4w�>V�!�)�K��ۂ�케I��F�B���e�(���]�� :��ro ���~~�
��x�v��G�[^����7�q]H�z�T"�ǋ��hJ��!c��ļ�1�Q�E�(����>S��[�¿��)]Gn ��q�ak�bF]�,E)S�6}h���s�0�	���78o��6����ܣfL,�G��� �)i������g�`Y_4֩�U�!l*�[J&?Qpv��IB˅�H�����+@��.^y#��$17�y��iQr��}w��Ǩ&yJAH�-����nR�ĸZ�a�"vK��=���=.&�$<�q�-���,N5*rt�m�촧g(����F��8���15a�'9��L��߁	�����gגD��py�3�3���+�60��V��\yY��[h�s%�˙����F�)>�I�Br�%B�č��.j!n�пg�rp������p��4�ۥh/��ʾ���~H���*���p��}��>	օa��������+בa��1A�S�,��g�}�[ۘ�s��'B��ȏ���@�b�Z�#�';y;��������4�����D`��L�R`6,�P��b�8?L��(�Tk�I�޷q�_��'W�k��p���S��fC����w�
A �.6hs8=>�����W����|*��L���b�k��U�JL]�oV�X��?M���.A6�>y�蝬�{�5(~�oȌ��Ւ��S�y�҆���a��ȱS�F/�=Ց�Ȃ�Uܩ±rYq$6���6_Tm��q��o�_I�sAhˁE��'ua�A�S%�%�Q���3�����r�A:�����r�'��dLE�l�לP�)�<߅
+����U�NsW�ⓞd�"�Gf����p��W�+��`�5�P��=*��#s !Y_~>����� V�	�!.�[Ն�w&1�PNz�4����\�u1,qT����Y긪E������({���+�M��}�k!��4'�C����������<�.����O�$�L|TmU��hԩ�ޭ6o�S��I)l_gW��H�w�;���(m,�vڟ���@I�	X����Zn��@U	�#+}�� �����׏�*�H&�/�sM:��8HA-��=��|��9�J����(Бc%�M?g��ļ�q/ʃ=#����M��M_��~Xl�+�ɮ�f������jD|Z�dWDu��H�1�Ě���9�Kn�W��G�0������/T�{K���wD������?� ��r4S
�CjS+9'X9�N��n�;�5����RQ8�;϶��q���ZP�\�h뼉L5�ռ�m�zI�7Å�s��gd��}?4S����J�߈����{,�0(su��+��K��:"нFDdQ��q�2Z�H3�<:%�QX��:{����=B*���bݴb�]I�ܘ�|>��g-[
�'u�	��>aTk����%?pXbz��ǟ�T�<I�['��7*�ӕ(����F?��C�Cu�����y7��?u#z>�@�F��>�6X��Թ���-6�L��	WJ�Ǟ�B�w�m(@���
@U�`��gd�<�
�mq1�#��d��%�4�gC^|@�y/�_%~M2�3On����%=
Q<w����6F:��J�;���pޒr���>ca�5̀۶��v��sJ�p8�aE�@5$�t�$�Y0ʿ��U� <������H*�y5�z�CEn�CH���=��W�	_���7rd��u	���EI�\��h!�5[M�6�Q��E��j��L�Rj�5 5����B��!Q��:f��yť��G�ŝ����Y8��6���1�>�<����46O������y&5����E�6���ݭ�yD�/!ezt�jO���l�������9Y6˄�:����o��iB�\�O�B���9�5o�Lo1C��|J��4yo7 Hz��c��ߑ�!ֺ/�p�%���vX�L(P�&�D�>e�{c�JU�uo��u��U�e�x�-�I�_�Ӎ���ˉM��%`��ѝl�!X��b���e^gQ�\���X��p	��a�5�ҿ�c���	���MG�dU��ܣ���ޛ\>}[C3�͐��C�{-+�w뺉3�eU3ñ �&n�lzV؛<�Ŷ�U�S��{�݂�x�%e5k�	���
���юm�̏6�K%�6��k ]D��t��7���eSi�xn�#��t.�ߜ>tW�VI���K�9xdLYwE{���<
@��6��8Hh-�ɺ=��W��Up��_���S�G؞���N7��ߜc>?�C���P<�^ي�=f}w MK��r#ٟ���y��*ӡ��h��S���X��D�&z�ʄ`��3�S�}�{Pr�w��q#&����M2��+�0d&�NZY��	���6g0~L���lD�BF��g=z��{�WiF���G��L����0�.���i5��d��gv�k����ܴ:t���nw]�G�� %a��^y%e�[�9�j̓�Ѥ�̗^ti��	�߃���L0Ƽ�&Q店�tX��������!��_�2+'U�J|�H&�Z/�cf�4��*�:�\wU��>�(.
�|���a#pi�.��\�ޫ�(��n��!qty\Ḵy���M�/흠�e��ɽ��lsH�<Ih�� /��&���~3�_Ȧ���[���E��%'�q	�"�EǺ��4�ot��kXB�1����S���_�;؊S7�s���f#��_(��Pa�#w�F���ҥ�����ѴW�G�N�$|&"_���Q�KhA�3��c�΢+Ud�]���*�?�*��T�M�톰h=�t3�h�#��#�^r��4B�l�e�((�pE9�V�0^0�Yߥ��Rm~(1�ç�~�-��Έm��$�x�u2�~��Ŏ$^˩��r����-K��� �ix�b��Űp�c�7	E#�im���D-�km�|ܞ%N�:g���znE�^â#7��g���7+�j�۫��i�����b⃷ݮ��?2�D-i���'�n1gn=�Z��AA�<IK�����(C��6�;gP�Iް�h�9Y:��{��G~vxٓ���[�h��p����N�������=�_L�!Z�_n�r���ʳI��2vC�������Jَ�7.Sb��T1GT�}��<1�i��mi;�!2�4pUTD�y3�R~y3�Ǎn4�=4�y*�t�<"wϪ��:+WN2`<*K��v������a,n����p��<%�n�;�K�)G����O��7A�X^o8�6�F���{1���b$���T�
���[�9L,|��gt��IZ�o1�m��l�,@A��'a�Pk�S/*�_�,X�������@?$ ���bc�6w�5�A0�'�?	��܋lBi�� �X���m��f��ؑ4S�
�&�B�zq
��΅ϣ��v�:�������H@"�Q�<����ػ��U}��+�w�T��2~��c��<���Pg��(��~Q�!�e��_m9���ԕR4N�g~�%KMi��&�I���a�P�jr��Ϧ6`���՛�u7Y�H�+n��V��٩��~<�y jv�Mb}��k���~._'���z���%V�m�[�̚���c{,�`PT��G3��B��A!q�l�Q)i��N��EjB��4�G��}�(�l,!)��ƪ�1��8�+>k�X��t���)�3&�x���l#�8O��x5t�ѩǽ�`�r�i�uz����y�YF�1�[�VrO��4L6����6�ɜ�+�4t��QQ���@�����gC�c8�X>���n�M�����l��H�y���1�˖�=9�`.��c����s�y:o-� ��ok_��;TBeu�~��9��Kɩ.�֯�aԤ�9i�j�\B�	���.���ڠ���oU��d�.��D�*K��7�65�Ϋ����9�jRPjq����� ����<����n��	����`�����N;�!R����b^�˱���~4�Q�&C?�L�̗�;޵�
)[��My��O!�ʽ$�j���3p�<6x����6/�H�n<X'��:'ǟ���ތ��"�0���R��i)ta��_�A�����6
"��Q!uV�"M3-�e�}s����-���Q�?�}���YD{���$�q���3�o�����K�9��X>�E�Y�t�P^�t=叉@uKL�{.d+�&�dL���A��>���Sh*��N3���J����ٖ�-��k����v���Z��v^[�&'5�V%#D��y�o�eR<Ru����Yec�er�b8�fP���V=����j��.j��S�jv�@㪱s�j�3��U⴯=ؐ�Q0�a��N:���A��M;�P2?�Q/ȕ��E�ϫ�������3ݐ�k���T �$�jx��\�t-����"3��u,ߧ��)X��շ�`+?�I2�N�� �)��3ήG�JGf�z,$!1�L�Ѭ�;U��K��,�Eu��ohν���4؛�4"X���o���m�`¼?��� S��}��桨of�$d8V�6p����?�09�e����d/�0<R&� V|GrL�s@Z���{�!����$=�`�=`F!�!�/3���YUw�^^"��� ��2����jz%�U�׻��bz�b��zEi2U���$�d5�11%.�1��`�=E�GN��1�ˮm��l��<��W C���Dbf^��'H��C��ɍ��L5l!�嚷��ﻕ�EL<(W�/��I|�����*g~<�����|�+2AB����J
��6:^8K�9bTzZ��w�Y�b�ʜ��RH�Y�h���������eM�
�-���	5��b�Og=3�i�#>�㊾�oE�Nb������M��.ϵ��Z�eI� '�m��u��7��e�9��w�f�h��F^������Ȫ9�q��$h�E��bp��w�B#7!�>!��K}9ON�A�%6B�W?@�K�mk|�56��2�3-��&���|�ӒK��<b]Wu9����Go��+�7Vqkw݋-m�89�&(���U{�_?���JD�~����UĎ0��`�~W2�2,L:����l;Y8�g�ELv1/��<�1�֤��0&=��l>�F�_� �dsCdL�2���x����Q���w&���Y��m2ҍ�7G�k|8���F{���3kh	A�_G=CLR��!�* /���Snz�%9�����plf�ER��N	#��Y��h�|�s/J�	m`E=��ֺ��)|3�{��@��	͞H(�l�g����
�Ľ+��7�����t�ɡ�+�C�Rh�u�^Q2��)%���(~�ҟ��X�iI\4U�}>�a:�n9��.���ƅ��O���
��/�:ub+��J�<�S�~G��a���a�Q�I S݁yb���5(�Y����Z���U7#2�4�+��b�sذ?f�R�^���.���"�gۦ�ʫ�g���c��9�U������g~����9─�����Iў�:����s�j�Ҁ�!K��ᦈ�L<t�]�;�W��
�O�2��c���&*Ġ�]�YՒy��E�R0�.X-�g�|���R����"�~��LX�x>܆u1 µg���F�X�z���n��_��?fS�K%�� ov<��{J�54��a��X_��#���D�h��^}�)O����j��I�f뜫$gR��u1��&�s����U5,�x�j��.v�~L���a?����*�J?2&\Ǹ�E�@C��K��Ѽ6j�4��ފJ�.sT����yDmF���tH#�&��ڇ�����p�ۙ*�Q�(n��` L��/o�1������eЀB�&!����Y�����"0Z��1�y�XU�Mj.(T L����X�� �q+��~����t��)�}�����+l_����7׏.���߀�h��I�5Ƿ$ۅ���Z��DG�+/p�s��"�-9���% e�*��`F���ꞟ�ѣ�e�叐�����-��ɣ	��_��t��. (R�"�T�}|(�YLN�W%f��3�e��^RҐ)����g�xδ��Љ��E�L������&�H�w@ �>ўO�p� ���>�F�?��{eǲT�4e�Z��S���C�=�=�έqX9�#�y�{�V��Bt�n�!K�� w$��X�u1P��%�GD����چu#�]�ބț�����m^"�0y�V�e�DQ�v��&M�I�լ)P�
h��������,OH�WM�蔏gz>�7��2Ϩ����ڛv�+�n��B�/{��?���ljN_RPěC4�~UgR�� <�)�pW�Q�r�Rw��쟴ڜPi�ԁh�|?�h�o8��%K�o�O�|g��!K<ZRr�j@�\p4����U��I�*ᐪ9�U���u���&�,����� �J�}��>8[�>Z�<Qj�2b��Id�i��^BJ)�%+u_�R��)&� LK�2-�����k���pB��1� ��k�V|qw��}��	�:�M��#]��p!�p��I1�Da[�x����F�t���m|��U���?���Lq�x�o�2d$e+F�9�� ��<��V���z�
/@2v��$|u�EȄPҪ�^	��t��yg�x���.�|�3g��b����<�U��C��K�I����m�3�����M�,ی�T��9��!	��C�
�p�L��X.&�=Q��]�����]�C�-p�,"=�ϔ�Y�$���9��
ȉI"�,H���s\@:�6ʓ�(�Bq�2&Cǎ��Q�2�C!N�˺b���1O�up���d:(W�9袶���E��k}C�|��1��m�p��~fhwէ%*��%Ү��P9��7��N8������ ��u� 0��z�;���I]�k�r��e\������ڶ���$(�l�~�C+P�����\�y�"6�:\�/�c�ܞ����QB�EE(��|#��X�{s8�����+NL��ҡ����]j��<�|}ڤ����U[��G��;�[3�h<��~��\�v��'�jpX�-A�Rܴ�T߾n�ۙ�هo�Ip�-"����sEΩ������ܓ-���'�Y ;d�>4ɮ�x�![�_>�}sT�-?P8�=�-�<|bR=y����#���RtV��+�O��{��Gt�z&33�4�^����<ރ�D;�b$��V���.��T �;<nBz���T���Z���p���х%����O>�z��{@�U륖<��c����%�����W��pP�ud܌l�n��,s�Eu�@��א��+�)ȵ���P���$�z&F����x�����~S�ܺ�� ���Sw��?b���B�-K2�)ْ!�x
�.5Z��-݉�S�E���|��5�ί4�hV�6�S�v冫�U�F&�
I��3i��!�Q6���܋s%�7�g�;A]Rd���]���}9W�{�a��b�f���h��FK���j
|�������F�vg��`x��5[��Z;��o�nW�n��OCOx�.B��H�5F��([}^��!�Y�.+������˲2�NΦ,|	���b���w�iEU��S�AaT2�M�'��~�8���ǩ���������	�g��n�oBO8��\��Ĵz�~���5��a"p��;����FÜ��?�\��z�I L��ue@R�5o���ly���V�UЄrC�h~[�=V�m�9���_�#��\�\@G��ޞ��?�Ā�H�yW|c�n���i�'%�c`���.��z�0�k�^�1�B\�P�C�D�6I��w��#|��5/ ��IL����-��r�ς�ϳS3s=�B�}���8���q�Ѿ�z�..0�����\t?���wb�fsK�a~�3IFL����Ow��*���S �NCD����i����z�D^;� �S���B���K�aך^��]c��'fϜ�08y��y�<�ܸS߀k�)Z��X[����z�N��9H��M.x����#r�cp��EMՒ;q�K��b/��E?|��{��b:�,�(?=�cŎm���×J�C�+�E�N�[��
l{r���&d!VYާ�T����Y�z����8�1VJ�m�� ��q�w�������'̒�i��|F�w3��g{��
A|Q~>�EִNG�Q�:��i��������rbٲ��&L�K�ͺ��������b�x$.��$�*���u6�8;}�y�|k�������k/U�����we��Y�V���j���u�^\�buR)U�l���M�T?�����u�E��-pR8���xy�xG��/�� �NI��Batk//#�_4.�D���i�n���m��Gd ��o=�UH����������IuC̀f7�fn�:�4�*MY�D�^�#��H�IZ�}'�S�p�:<�៵����S�8���|sZim��~�T+8��;�7�&�୭���� �<�v7��m�$҆n�����<{�+m��t��E�4O����i&�Lko�k}L���ʉ��B3�'ާ�?A\jgn���4�C��lH6::S�0��(���Ü.
Ǝ��9��	L�ٸ���w�s��y�8�*i���Շ�����;h�a�ml{xiNQ��4 ����3�:��Gu�p}�&gxA�E��?3��0��l�UEP�R	��b�̀���\6'^j��/���X��[�g9��Y�%�7̭�f�9H���
�~�ǅ��Gt��=*�^O��	�<{��2>���p||u�s<h1�}���*n�l�U���H=`��)O`m紉[�o�x��?��4���0����\�(�-r�R�s\�Z��'��"�<�7��G�w��>�X��\̆��D0豀�0��QA����ow����j�Kj��:����5��S+�qOlr����Z3+v1���1T}��ؽ�{c���b5���k�����%�5c�.M7F�֠w�D��b�|T��p�X�%ڴȲ`�p�Sw��Q_WH��N�ZA�p^څ%�,c���z�ZG���������f�>��*�m�Υ��?Mgc��/`X���ڛ���ͽp�VT���6��ϡ��U�rF҈"Q"t��t��uάī�g����
y�,%uwh�ɽ���#�(���\��S�]�|��F��}�J2��K����F�ry�a�#>�a2h��W	N3,1���I��Oa�g:��d�'�M@
j=�d?��T������^5�,��-�q������YbWTǅ�b^/�|:���2L��K,�4i<�s-�:�{
-|�O�)mE�c�a ���e㚮/b]F�mB%�r �Pk@��Y<��3� ��>;�1k@���y�)�YӼ�k�Q�ɘ�E�)׾�w?�:-���HlU�p!�Z�2W��V�,�d��S�&�S���rY��Y�
n�^L��DS�>n1oZ/��U��qK8U�rm �h�6Cݏ���;g�E���L�d�ϭ> �V�`	�c����E��l�F�"�3��Y�|�� ��UE
ibbq��w�#�^�B[�TQ��)�?�Vz�4Ʃ��^��:W��D�9a�Q,.a�h�5�����n�7���e/1�[�1S�Mg�|��՘�ո4�h��9�)�jl���!hsj�n?�2�*kK.4;�ԝ�_)h^�}��ʏ!{:}�R�ɡ��:�R�ȡ1w�y-5��7���7����HkCY8��k����<�#F��!�#G>μ%>�7<Wջ0/��`e�N6�X��'"�Vd{�@7�My_��C:�-6�M1��R0�Wץ|XQ�[}�؄�1��� C0G���^#jN7���6�"/��(G�W��
/�c�40��E�<
��b���ɥ�u<v�jb�D��}|Y�P��,�8�$�ʋlW|3����]{_���!:�c�%��qZs[Mݵ��8�V�N��-yt��fP���1T�������)E���ȋaZ���s�¤<���5Z/�Q�Pe����>�P�}�\��Dӥ�X�sH��Q�p����E���k�K���_�#��]jU����ց��;�XG��� ��QZ�L��� ���q�lf;�҈
�E��4r�2���A*�;-�O�<jSW�Hb\ޢ�x��fHt�KM�.<�ǱC2:a8�i�x3�I�pI��8]ĝE���m!K&���/	�;�O��{Q%
�w#����T� �}��_P��D:ʠ��,�$`
��>g��]�J�X`�H�?��7o��@��������hc{!\��_{�i��K���e:v�������Y�D�&� I�96�����)(��\� d��w6�m0֎��ـ2h��IS�Z�@t���������������oV��|���"]�i�5u,�� ��U�o�����~�DLx�?��ց��R-RH��늹�%YUm�I3��˸Y��6S�
��(m�j�e�C���^>��,���r��qr�.�_�("*�rEN�7}EU�C{�|W:��`�OՓX�7���}d�-W�tc#���>�i��sN����|;{���@�,-!ȖJ�B�e"7$\?�i`m"��6z��i��՞ G���q�߾_������:��h��E�����|A��C9)�g���ɠ*r��|/;�nӃr�k��M��ᨯ1��T�-U��ˎv���47��[�0�PH1X>�b����;��$���i\�3��,'��:|�Д7��z��-�,U�u���0U=��
�Z1��y��F8�7��L��j�˙��N��@�섑;����u$�t���a6 ު?����ԑk앝��8����^-��:��9U��?��؀$�z�T��!].dd��pcC\fH�����%�!�L���l&�9?�T��Yul.�S�ܬ�ݱ* %�({8��Y�F��PoPf��X����3���+���R���_�A�W�)�|��an�X��%ٹ1�xw�ݵ\+w	,	�����8����DSd{�k����v�ޡL5�������2�)��iُ�B��Uo��1�Vc���%�P�XC�Ywm�qR��eo��v�J1f�sɃ9Q��� �BJżE&��tc��&�/q��a��\j^[�IH���j�:$�^�e��g��<��$u�#��hR��������ɰW��֐���Z��֍��5]�5d�QvBxg���?ugו�9�F��>D������4%�;߶�E�V��Y��E�"��^$�8�
̂>G(G�o�q:���;�՟υ�E8j7﹤����R��z<��i��C{��<����`s0������Hu�e<�\�c`�	�>4��5�,s�;�h;E��'Ѕ7<�!��K�$xT�����UʰA��M-1~���hV����G��g"&x;��dΞ���4�b����<F�ࢵ��qV���&?T3���6}����p�G�.�k���S-G�A6��5.m��{L��:��,�������'*��~;�o��u�Rb��2���M�z�(>#�Q�|��"�/ډ���)��H���|9��nB�UɡeCTn�5Q�1s��&\�(.�7w�cY�yu����	��&g^œب,[�V8��hU:Y�nDg�·O��x|�����n�<�u=�+f줛E,r���l�@&d�)��/�9&���c�P��_�͙��V�I�& ���gDL��<�J�Mk��NwR��[�GE����s�[��J�����9�d�gU4RfM�r�1�fZ&���]b��Q�Jhh,�z�����HǼg�R���?�����۱�P^T|��w��*	/<PO�
���<|be��c�N���]<�RW���쪬{�)tO+����LA�^�����$fy�f�y��_�5=R�?�u65�.}�b�}	�uwTXn?I|0[���*9̭��o[>�-�
����)|P���\��xne5��U��tr�"����2~���⸔+K��i-%4��Sc+E#���%� ���B�._`�ql�lw���:�(�$~�CJ.�aQ!����QH���M��
�%���J���[zs!����-|Ql����J� ʺx�ަ-WQA�t��d'����.3()§���4XH�N=��"�*�=�=&�x�CM�?�WbPuh�	"���F����(u_�L/t~���|!r v��>��GX��bY�*��I���`&	����`�ZmcV�qk
����jrFH���'��Vέ4V1����x���x�2�يH�����3?C��#�~���:��9�j������$�����ŏ�E�ʙ/(�6�ց�|Y&��΅��5�%�q�*��nXi�?�L�y �x:�;f�Al�FZ"�q�RA��#x�����u��M��nk��r8�4��`��Y�y]�X0L��P�ΰ2����'��&�sH�j��̃��۪����k�k�J�@��$����ik|E�O�-� r�KE�6�=�6�ک�%v}:395�_�e��+e^���jG��}",j�h�7�.��^Q}aQ��#,:�u4eZ�e3Iɤ�`O�s�=� �J��|��������<��p�1ZS�a`+஺��5��V�&?jJ�\n�]�e������ؑ1�r�BZ�����">�˲�v�D[o�������h=~_��i�Rz���*�����D�¶�z�b�V肏˙��u�	�@d���
6B Ϗ6ߑ��)���)el&���ÒS�1�KyKŠ�E`��l�D������wy�U;`������@#d)��=�QΚgy��i��CNW�1�0�N5��4���UfD�k������T� ���3G�yL
���ĬZ
Լ��ӿ�=B��b�p��1�^k���Eq+��t�ny�*d� �ѣ��9�����mg��;Z�p}W�f �<ԃ���mn��oA����2���%��`�K�)]�WQ��+t�2�T=�:h�fǶ�4�jJ@����rm�-# �h���+�tE���bd�	�mʜ����1|Ïb/�����2���b�!}������7E������9ŀ5Kw�/Э(�^p��@�f��.�Z �{������h�LU;�Kc��K��0�Ȯ@� �n�Cs��G^���S���xn��Zż�� O�)�Y��w�e�U�4i�ީ���4E���;�v*A�*l}�	4�x-���c�t?tf���½
(MNw��}��KS�g�\�ԇ�8h���M9��8}�����j�"9}g���7��~��Ú /(+;M`g<l�fHBf�ds���ѷ�F��n���fp!��Q8/����/��f�T�����py��G��i��S�D[�������c�Ĝ
Jf�H5J}�f� �����s���(6�c~��2���9,f+��Y�'��{�d��M(iA;�	��qgZ���9"9w*JU��h!�w���^��f�fj�*����T�?|��A�<⑇f2��d��ɚG�:?)k��i(��� �'3z��������U6��+���Y۬gʽ7�k��Æsػ˻X��Q��/�k�=4��V�g���V�*��
<�4.%.n����2y��·�K���f��_�r�m��y����b��'�pj���������P*-��@Ìw�ԅe�@3���_�h'|��w���5G8u�.�í�/0틆���4�r�A�H�ho^�K����Av����d���J���ݪL��l���+U7��'�J[S5������j��p��m��@֘�cBf!��_�+�jS�Ez5���'�Yl��v����
y���)*,�И�����BV�d�ڵ(^��*���E����v=�:!9?��̣ ���z�y��Kgm����BZ��B�T��vb�s�S�Q��j�����)3����J����g��,���#~���.[E���c7�_�C�؍��lc:����������TV3�P'T'^cK�0�lk]b�C�|p�L�%�6a�5VOҟbH'�SM��N���(,�/�#A(�W�5��
b�%b���e���4L�%[~c�� Ƽ��W_���U�k �P~"EDn�<:��
��	����`�ڕ�3S�"e��ػ�s�7����X;����P����^tX�AeDg���J�g�_Ʉ��X7�8j���H��N	yl�קAp��Zڋ�%�_,�|�>��y��F�=��%j,���ђ1�o�u��?wA�6U��s�d�����_຋Ĳ��+���K���Wtm� �.X):1^�k1!�6�L���	�ek������M�q�q�m|׉��9�1ud'<������*�#���1���� 7�ZQ�F ��>pߏ	l���7�r��p�}^�V�ڏ �1|C�5�'��E�']t���4�u"�G�즅�aeԝ9<4�[J>�Eכ7�pJ���9�v���&X{4�xJ/�0��-�{R����3 	VE��u��؋�Ճ� w�*��[�Spճ^��Ւ��|��\[JM�Z5��	*.�ً��V���H���5�����ĳHmb��i�{�J4a ΰprݎ�V�h�wN��w��i����R�Xo����I�۴+�-��.��[&�s��#C�9Cݟa�k��=�V3�]�2&��<�ʤ�Mr�~��@�4oE���b��E!�_o�0�1�~�G##����oٺ[�kQ�7<Ǳ�ra�Z�������(�L�Xvք�����g�����7�{:��0��#�b@)pY���S�G�p�Bs�&8�T�u���r�]?;A��Գ���*��Md�˰��>ｙ�����m'���8��_ͫp�� � ����}vV��F�͎5y�����.ߐB�N�����Z�C�g6o�>(��XJ{z]Yj�J!��Ϻ���u�������V�DR'�Q�@�~t��?cΏ�����Ϻ�D�����Q�o�At�F��`����>A4}�]��Ha��T-&������]UK�$eY�Ǘa��1�_���Xu�k��m�D϶S5;!1�#�Wz��m�$;f�����z�>� ��a��S�N}ق۹q���Ò_�t�/��G�1�漷"~z��D*���2�ָ�`��ս?v�t���mXnN�����dw�|�[���� �'�3WJ#W�VƋ��^�c0��*U�G�<����*�N�D��lp�V�#�<T=��ml�+�"���`6y:o0_M5�L	�2�M�S��-]�����/��=P�C7;Q7�ܪ?a���
CBb��v�+�:��;����v������������������pOB.�t_�ޣ�T�!�§t@�<eڲB�۔7��{5��w<�	ԧ�J��Ì�!�A
긍��ٙ���.�Ԙu�evŲ�x:'���ffgr:N��|���5W<KBy(�&L>�����.���sl�x�o�[���]�
�W��1�D���)��ub�1H�55��&K��ye��4,�=�>�5���[�<S�֩��q�!�u|��&x���e�#'u�6�mj�8�5~�p� f�A����<>!~:����@[K��1��(���	,��j�_�n�dm���y+�K檕����������s�ɭ���M&���+"�~cƛ��x�|o����j��(ع=|z�4�QT�&.c��.�Ms�"�����)~�q���L�Chg#���#.T�?�0:*�~l2�'gp���?p�JJ���Wͻ�2b��bJ�eb��#/ct�j�X+`��4�.�nϦu>&���o��~Tr�o�pf	��k�s���s�E��B�M��K.(����Ņ�������~2$��L齶��b^oo���2�0��u٩��!k%�-�]$M-�jn+F�7D��՗-��d�}���b�Ap���1<��RruXkJ��uV�I��\�8X�Uțh߬�y����i��mŠ=�(�Q�A/_�����%��L�P[�U\��9I+���v�=�*b���?,'��\N�>�q�u߿�0W%O��Aa ��f0\|�∊�έ7�b�,����Ǧ_���Q8\N�~C����6��bP����t���W��~Ӽ�ǀdi% f��D������W{��ĘD��I��p��e�����p��X����j��D�J�������m��PT�M[h;�_7H��84�'8��9-0����x�:j�N�F��A��_`��ô����?1= Sp0?�¥����X��F�7� A�T�䛖���	85�-�"�M;�^�k@H �rL=�g�ŀ�,,�KF<�umʯ9�wE���#3����U�;�"rM���.�K�I�e�Q���J#6u���#Я���yA����c��e`�t2��� �[b������A�T!�qt!d�d�����ĳ�[h�6,,�A�&M��a/²���R�ɯ����,&��19Q���@[�X�>�^5�ݶƆ�1��wC�9��7Iz(�޻��d�%��{�I�Ձ��!;����(���<�>��U��>ݼ��ئ �^�А'-�z^��^��H5,�Df@�QL��XB��䖸�OU(��Bm��{d��-��I��nf��iz���-ۤ���*+�2
�d(AK�U��O	�H�0_""�W��b?߯�3=�$����az"��y�/A���A�jP��2|8�i^�&����!&�g�բ����ˢu+�;8�hu�}c�"������ք?�or�A<�bF)�u|�c�����������RKEWA���t����3���älrp�D$�2�y����
5�v5['z�����niΛ�|�y-�o]��G2��l��*�	=�/u+D�>hZ��90I�1�f�`�
"�0�37���>SJN����F�)���UΥ��@�̳V�2(6l��ˬ)y��{`����� �� wh�p\��ߢ-t�+���c���"�^�e�g_(�<�џ_}e#�ٹ����S��J�#n����]&T1��n=$`fXu����<��`�<��G�'\�;nP���ū���{�@�p+{��obrǠB�K�,<��4��]4�f���>��3�k��wt���?�ŎTñ�ѬjOq���������I�Z'6��5�5�����2X�]t?�s�
={������O�I��CƆd�28s�0�G"��~5΢_�G�G��������zG��RɁ����%����p�a�2-�JW^.?�q�
o#�$����ﴋ+�<�����7�O���A��&#g�ČtQn&`4�ڻp��_���IN�iR�\	�$%�Yz�|p���LP%
x=5)�J�U4��C��:D�]�nV�a`�裫,"v�z�g�Lb�V����2_�} ����#�-����)x�3�0�M,;!�m[;ݣ�]Jj>Z������,���Ҏ?�V��m���g�����[J��h�{�;,��@M�	�^ڊ ��Аnp~b��ha�]�pm�YՐHs��[���Ȟ3���h��u�'\�����?���������jI�H�wS�C-�����Ϩ�s�
�Ye��ύ���<��ZsO%�tќ�x�A�� �K�*�}7�^���eğP*w5��D�F;���h�˃g�����B+*�
�F� �šR� -Qr+�^�Q�AB
�߿�e�pL"Y���ı�p��A�w.x���+����i��-�:��f�{Dp��`�X���@O�b����n���#C���WG���PY ��sT@B����N�u�R�A�n;Nb%x� &;(����$�=kg���E;�54��`A�����U�ո m
���"o��8l�+tD����>-H h�d�\��L�-Cћ(N��>H�j\��|i�CD�O�|oX�1',�fp�����DvJ͗c��)�څ��]ˇe��ЃF�%�RT$٘�Z�0��5�UƦ�(����]q,K����t�Y�Y�:Ӫ������D�8��tqSBMy��5�\�;�\��X�.�0�Dٌޔ'�1즣jL.v}K&�c�:j�+�bhE%J�_����W"ZO�7Ȟn4�\�=u2*��E�'�z��'g+R=`�9�z�K�p%>�xr�? E��,L�_Az����H}wl;Z��
�� c�G�ު�o� 2b���:��6v�	òD�?(O�O��|��y�6��8�/�b����8�����2���6uW��{бf&��`#j�����YU_i�W��<��:Δ��5yN{��k�YA��N\D�lzr��
��z�h�Cm�)�?'[��)~�C��� z�Q���?B�kW�a���^�h�V*��F��\t�&.���$7���v�1���>��lm�l#�]��X67�}P�V�V�2���ipi��
=�+���P��-��D��ei��+3�B��I�H����Q�(9z)��*V?�y���A�Yj#��)Όug齹�aKҶ�S��AA�Ȑ�ƌH�S#5P|� �S^�;�"Ak%�>��?�����R����7HǊ;�13۬��;}�ݶ>�P�W�s̪eCL���������M�x�{�l��[��u���l2�����>�������"� Ҕ+���iV�>�tӅ��Y��C0;J�҆E*AV!�5n=�9k͞�!"u�����b�Ac���|�4#*\�r�qSۧ#��M�V��U����d�'�8x�)*ӄT�*p2&�/�,�w�"��z����s 3+ك�2��y���BU�V顀<�0�gm�*#ޕ�-�L�>b���	}	���ɣ�C�#�R��8\�,��6�g�����)*�!�G��`|s��5����G�<��%���w�=�,�	��G��=y�h�a�ծ.��HL�q���Sv�ZX��dow*1ۻt�#�G�[!�<��0�
��<	���0�H�zC����T�,�����z�w/�A?�U޳��
fH0}vףU���mXa�\=�47:gN�s<�DGt	�(I�J��	��5�2�=Qm��?��2�%�B��&�ڗӀ)@4MIid=W��Y��N��`5 �%R ���C���"P����`���):���fJ~;���:���)�!���[�*��]k�rx5u��W�օ����s��v�˳N�'ڙI��vP��=��ϔN/����b�����#�ۇvO��cr<z�*�kqjeRf����l�_�G���$���\Tn�>4ӊ�iq���\���" S���Tu�2�������.����N�A���$����ƻ�O�٫o_}r�E:�P=�M?�I�L%���8*�ea�O�(JV,r>M����q��=�$ʎNl>��*R����ؽ�=(,1�����T�U���.��X	��c�˫Rd0pK6�Rc쉄�sJxؙ� �-r�@���`RC"�<"9J˳���覤��fA�k!�mM�a��f�5���$}�j�>�sm��!S�S�/�R[��:ő���>/���p@�g��9�[|T�:Xvב���b��M�,{�`1�-8�Z�z��c\�J]���ȧ�����kZ�z�DE������'�%('�M���`�	��8gdIa�g��ƆQ �,��0��J^����8��WM������z�2:���f��/j_�wwL~Qr�mn/J�Ip\��@��Ç��+���*�����,�2cݦ\
���,�����H!Q����/K6zQI��w��O��f|g��8����E�c��ʁ��� �{�V�{�����gC��F�2�I�3�0�2�	b%C1��{{��?���>;��`�� ����z-��8�t��L�ȅ��ns�U����vi@�r?to�c�	�~T�R��11����w=������"'�\1�h\�|u�1[��r_!Q3�X��s�(zK��@�0q�u�}9׎Q�y���دB6L?Ud4�X��X�k� ���d�4(��fʞ�B�ݡO=�s8�d�)�0�!�FeK{yt�`ǋ�|���9bצ��4gs�8.�1?5���?��!��.n�X�5�Y#@�Q=���B�� �\_�*׺��Td(�6�c�*Q�-���ȾZFGT��ð|���7�nt%�N�gu~¼f�V|f��pmSN'$i�|�v�n�w_]x}�.6� Ň\��H�	[�գ�lN�qBk�0̻	9��ʞe�X,cجy�Y7�J�����~'k����w\��9�@˙Q\�T�R�0��l�㩙�ys߳�K�Ғ���/ !mg5��ɖQ��W�4V	�>6�#���v��	��-�QI�hM���{�h����v����$�AM����⦃|pﶺ��M���Y�����3���D4����tZ��U0���:�O�ߚ�!&��'�!?^3�o�,-�ʑ^�e]�b�`�(8�a]�|:	�`�F��ݗrX��[�RJ�
&��=�@�;>Ӎ$;}�-;3�̓��S�ao����mK䚗�b�hQ�)O�zY��哓��/���cC����x��`�)a���F��(��ɖ���Ą�
��_-5�j�����E�0y��M�T�*&���"F8�ʻqF�~#!F����zF���d�zGj���j��3�!y�{��vB���P����Gc���\K)�h-^��� ��nzY�6]h���L?�U�[H�M�L�k4�V������D�q�kk�^}&�b��Ů�՞wQS���I��h�����K�X�x��y�S�b��eb�}�N�:.9Gd8���.�4�k9��|�*�٨�Яz��y&$���m�|M�3�TI�W8�[0�Ի�tgR�m� �c̷>\�*p&��p�-FG�Y���z�wn��nh�������Q�W�P�5�Y�k{�X�������$Дm���S�s 'ʭ��@����+p��	c�f�����lю�~��_��� �f�V4�ϟ��ǵr��`���~�+���ץ�ƙ_����y����gի��u1J���J)�;��5���o�o�>�jg��V�,/�0�>}�Z�o��`��N��b:-+¡���u��Ĵ����1�u�Z���V/��\WTe��Iu��D̬	sR���#���y��t�	���)f���
1���#�+��q-d�Fށ�a���� (bl�.D�a������{g�q�uX�ʫ֯�~��?�f�4��@
\ U;*Y�+��!5���k"|��q�,��J�o|��NPi��뾁�� �*���*3:��ß8��12D�Y��1{	�;��/lX�1L��.`pV�s��v�|��!)��v2hX�jg$�@����`-�-F��mF���ǫ�4�]e�=�y�Ř��}ݓ� g�"��rp�Msf���a�y�r� 8� ��K,�]�$Q����-Mz���
ބ����۠B�^�GbBC��E5��J3#������YեTr�_6�M�q7��v��#���$tvo�� ����;\`}���;��k�[ �W�;�&Z�n�K��h7%�����|���b��uIw����"�������=Q��v6��}���c���Q�BǕ�`�k_�����jD�����̉����uS?	C�"U�1Ƴ:��h�U#&A'i�t�A����o8�i֪�׏W��ɹcP�\Ъni�G�*��0Rf[���F��ܿO�bٷ.�~��5�w޾��٬����`-q"%)o-"�WF���# 6��8�ש�VO���|0�O�T��P�I��Aݜ���|6c{#F�#�#�3��Q�@d��� a٤i��M�ړ�ݺ ���#d�|��9,�����*[�(��7T��,GY\��6I.�N�O�f�Ѡ�+���JK%�g�ʽ�1�{\���^��aH�l�zN�<J�у?x��G笋R��p�h��,�7m&F�J��8&z3X�r��SDY�YA��t�w����Z�\]��ʽA$�+K�k�e��Ck�Z���,ӷ�=Q��6�d��8����߈�#��\S�m��m��~�,,���؁9wl�)f��<&Vm?�'U4���ۊ�2��-�7ӌ�	�YXu�=j�>��հ�b�{�.'�}p�<2!���*>�
A�,�/���.�40�"�i�X�y����-�D��`b�z���� �K��O�����_��D�/)k)\yH�▵����]�ė� ��K��.K�۷/©�+�H(����6.��2v:��~z��Ψ���yP��ѷ�O�<��R�ź�ٺ���@�t�8cm��Ao�H8�̹6� �y��h�
��K6�8���jx�Y�F�-'C��5��jD��|E<��E����o.��Y�Z��گ?�D��p�6�������V@���yi�Z���ٽ�6���ٰ�Ct���+ɂe�t�PO�Y� ��Ce�������k�_�?5*D�]a8jP����R�"n�ʼv�L=�1a�s>��D�S�8��.�D_S�]3bR�����z6c2���V��	�;[t�J$]��k긦�?��_���f���7�*s4v�.0$0�m	���{>'(�(�明b�Y�E�a���� ��G"o��&+
o�i�^�]��_���P�V���w����� ]8#%�%t��1����/P3X-�	9CI�X���3'����[��k,�Z%/��L��uOl��9���O�A�K�����S8q[�+:��Q	��pC9M
�(���ޢ�P�Ɗ��.]���"f{�V��A����AE^��|n�&�m!e@�v���9������ߕ{������;� �4_2�*|ġaU�t"��mٚ�a}���!SY�FE�F�w�\w��>�0W~�pA+~wo<��G;��}�H���t��tg(&z>4C��R���ǈ��X��-���
H�9*�)�fw��b�\Y��t�����Q�B��{O�o�ol8x����H�P�5+Vč|�fFnc���h^�C��p�*�x�"�=�X1D5R<�F��a�)+���b8BVsL~�$���g����U�O�
T��}͐����O���t�����1��]5C#]1�Љ/����,�Y20d���멧[�4t�b��K��,�`2@
{�q����h0`m�x�m��G��0�i���Oqu��𸎸ԦC|q~M�������O��h�f�g����E���N����a�!F�נ1�+��4+Y�;#޹���@w�װ$��!��F�����'��`�o�<|v�DobMw�?;�6<�R�����#���g�9�w�rV<E4P��M�}�:����_W
Y�Iw0�fW@�~�%Ș���ۻ�dE���'��Tl��P���ED� �M���c)�B�5��9�Q��4O})Um�(q�x���LрD�EG��Ӑ���8I������.5J{�b7� �hUF��e��> N��%���� ��l�ٻ�/D��ɗ�i�D�q��u\0��'��E�h�h���)/%t�p�1��\�����;���xG�q݌cn�-@���n�3��;1�r�̉�.�h*tW�k��xuj�,�\9s�:�G��'C����)�$��p�쟘�|�/�acL��M�;���[��Pe*C� j͍[�@�o�xGz�^k�bI�U����	�@W��xf�dN���� �:�H՘P-|CV����ذC�n{8��c�sOONf�mx
"5��;�uG6n+C6Q;񅳸��˗���u63��q�����BwG-��bǹ�qq;��uB��k[��^"�Z�U�V��챏kb�i�X5G5��������Ab���4(�,��K�l�	����]GG�f��4����EЌ��)t⸋fD��۴�`��9���ޖ�O����М���pr���lep�� 8Y�$h����8B[���		-������"ipa-�\z�y����솈��?�L/!���o������(�:�=��Q�1|ƕ��wA��i�Vy�;��ay@Uџ�F��\i]?�y6��.�� S_5\��#23��h��4l�
��^�'��X�Ӫ�,�7њU t�{=3FdͅL�ݿ�-� �e�R����>�Y�L��e��a���a4���v�QC������6i=�^ݫ֑��~��%O���yR��4b��r9�猔��~���?���HVyT��O�)�Vc��a�%`3�O����W��نM/�M�L��$.��y��e]�C�+QϭIϥ&�Z[�$?�A��5cb�;��tZ.�}��� T-/B�+��` z)�ߋ��v����B��N���Q;�g�����?��%�LJb�;>�"h�=qL+(S��D%r%���$�O,dC���QHb�-���ܓ`Ċ@iT�J���K���fMt�cT�-�r�/[4 �_�/�U+�0I�Ҥ�+X��鸇�\I:����_��g���*��1���M���k>��M=0��\k��p/,_Z�B���_����g����BU�(9��4kk2��^��1P�Q�T�{Z�<�f��q�Vr����&��[n&���i�A��3���;���4�X�\k`"��#ԍ�Zx ���+��>�ø'�5����6�2RY���NC���v����Q~�b���]��^��hS���/��o/r�T0�JwCE�����~p��tn �o�&e���$�>0ۂ)���:˱����{�M�)ܥV��4	��ߑ5%��[Q�xmX�Dr�F��H�kZbP�#�?�Z�*�&�����Z��˰���&�t�Ro:d�E0�j�u���V!e���-Q��%�\��qmnK���z�8�|e$-��3X?L����*ѭ]5X�þl,���s{��a2�\�+�"�Qq"@|3p#P#�A���~�}�>Y�0�ko�٨��D��Ƿ@�C�5�\�tnj�%ԳY8Vx?����-[H��U���d׮��h�'G�5������ŧ�'딵��=y��� d�%b$�o�F����S�|4((���Ƒ�3�-�"�9D�
ʏK�y�O^@dIf���>��~K�u��(Q�ܴ|ҷؐ�������
��Wn��Б�ބh���+��5��S�}���嗱o�vf|�Ӽ���7�,��{"����vh U$`|_�j�u�!��nq���J�+ �:;y;�\i�bN����t�+��~����,���0F�VΔ��Q���)4P�o�Ɨ%����">��=z�����bϿ_	ʣЌ�#İ�"�<�&�5�zI���u>�Au�Mi�
0��N0�^5�(_S9����C�G�ص�|���⟪gn��b�2D��J�W=���Z+���z	���`W_\<$����9�M�-�e5�	�%�Z��!�j��4���J�	�M?�����W}�ư'�����Q��b��$����\v�#��3i �8����l���HE�~�q]VP$V��	�p�����*m�b`�P>_��c R�R����?������׸�eʋߺ.`��Y��d6ަ��}u���,I��ST��hc{p�sm�10=a��l ��F��<����C�2�S$PKf��>�VH�_��M�!�y�'�w��W)st�Z�,qoCe�å?W���Z�aTY����[������hO ��]�R��A�d�GO�;S�;���˦[2����<��ܞh0��}�/�״�Z��*�W�/%+��p�ɺ�޹;B����Դ�8
U���v;�vR�}�˲�Tb5!����C��m"@���t�g˝�L+���PY-�1��ze5_3�5����S͖�Hms�a���'�Y� ���p��ϣn�:���]����`?j���W45޶]�Ž��@�\���O)���Eѳ�&v�
���h��f�n~��hqM�����o��Ϲ��OE�¾B��mQ�+7m�T)[b�I|��-��aN]���a�=�H���^pB�~S�CCA�3;�{Ɛ�KR��-qŠ����de�������M�u��°H|w�l,�8��������y��(��3�&��AILڣ�u�jA��W���4��񮺘e+��Ǳ"�	�C��Y�}rr���E�7���(�]��G�~mi-�����o������N�%T���%d+�ܓ"�N� ����+��,� ����r�d�c�~mZg�9�0�+���A���)�i/pq�i h�ɩp]R����舢?��^�%!tv��&�#�?�+
�\�[�e��k̔�����r[Vx�,vﺔ���W��S������e�ޅ�=������6��!�^���fA��
��Y�[A3;Kv4�{�G<"��`ZK/J��KfG3˩o�VM��v ��AKJ 41��7V+���59�.�=��$�L�We���2���8�e��`�}�|�"S�I�V^ٕ�Fy��8�Py��/8�)Ә��	!����u~�DC��Sv���?��D���̲"Q��}�2�_M�'��zC���r��:*�Q#]�zU|S_ c
ؒE�[)�C�ʾH� �CL�13�h���tR?��n�7�}�����Z݃����d[��P����}.�}&�ͮ�
�J��� \0=H�x�uM�
V�����w
��!-�}��7��1K/�!<D�ܫu!�ґ�PPsc>	sٮ�Nh��Κ9r{4����ݷ�u��v_���hB��>0Ԓ�Q���׭����[��ȑn��� 	�x+3�	��u�}����:�a�Y�T: ���yI���:Xg\��[��L����7����j\7,��5�tt�SI��,��o4�i����.��hla�1$Fu�bM�~?���(=ot��}�(�2z���4/�z�H�XH���o�r�k���	�� )�p�l�ӈ�fU�+�>Y\١dX�Q_��+�ͨX��fķ<D�C� �^�@_Gwn��Eu���U�(���K-�lZ3 �<�"ed��lJJ}|��B�ˮ+"H���S�D��N5�Cd��	Ld�
��z��'*kx�����I���z7���G푶tׅJ1���i�i�4��,�}3�3�%J����u�ѩB�-ʗ��O$7c}@����]|�A�0Y�ؐ�H��p�G�p��M_���{�A�]c���F��W��5ʺ|���J��O��6����M����f��[���Ř���	� ��Ҡ�u�]ͷ��t"	LD���^E� p��y�S8�j@4�w�;�ɝ,XJ�?l@|$�}Cə�����˂�M�\D���s:<�PG�I,�\���и������X�F��ڵ���sz|)g�8lOT%C(o$b{�%`<�|*��O|���Ơ�^	�Vi�Pg��T[wڌ�m8��V}^ָa��&~�#5K�ڀ�>������O��.L��6���$%��p�� �()9�P��ۀ��O�@���W�p��AJH��,?�P-)Ձ� ��㡅�;O�(�T�I�A)��,B F~���9Й�[t
�9�n����o���q5���j�r�:�Bwb����e~{��mC���qg�\���>#*�ҋթ�-%�\^6��»a0��n���>��p*�b���{f#�:՗$�t{%����]��T8��WkљȲ$R��5E��;xu����wTf��U����mu_���^+��i�@P�Դ��w6 D���'2h��L+4�/�v��K�D��Ԋ���"������O��6�5.��K�����3�,��t��<G��nI�cz��u0z��tjR��ll��GI]�!�̥K�� fe�r,m������x�a)��ޮm�&F@5(�g'L�ln/����y��U�ˏ��پF�u�׾Aр�1@*A���d���e��c━t���d1-o:��<0يN����)!-a�j9���=� |��{A)�o�,��aI��LOg����3z���ŭ�/HV����Y�Vb�x��X�peF�E�����yA��'�� [��&��w%<�@��ߧ\Xh���/<�[��.4��*xU&|�Z�;���;��7��"������zDm�N�u�̂�N�?2�G~�t?1�#�H�&�./,;g!H"Hd��d��l�5����;����ח�i��c?�4�[��-�Tb�ấ��ť�&gl�O�f��V�}m,Πr���U��> ͖X�/�����@R9�/o:���7G�h�8o]nѓd�4��q3�|��3�}!_��I�X�W���t�Ֆ�,����1�c�NR�����eY�	��s2�:�笪�K/I-�'�	�L�\"�	�!��~٫��z�<�e�{�������B�6,տ���47dh� �<�;�;X����$2��������3���`�B����\�%Cm�x��7o���T����2�7n���z��ou�� $x|�R|�>δ���r��h[��c�t%���yIq�t��{Zu�+pSv��K9�3���ܫ���s��D�>Y����I�] 9}>z6���n��\�؋�OV}�Π�:\��\9R���g��g�4[�wF�	��W������ep����O���W������~�Xy��4���Y�2�E; �4��J'�vD���U@EW$��U9�x�TN)�!z�~/��p�[�YN�F)Z[_+|b�C�x����AK��j;��-�����?;��r�w8(;36��˝42o�J^���Gތ��3У���1ꈄ i]�ɟ]�O���Ǔ��'�RRu��o!3�m�k�t%*o*ʩh���]7(-܉��;�ܗ?�A��dطǤ�T�"��~���JB�
�� ��O&Yn^Ǘ}�Oa���ؐƋqUɌ1�0����<5��&2�iiuR#[!9��zQDL��g��S�-���P�q�5�
����T��'�;�DA��M®	�T0X�q�'���&�~-԰����R-쓞��)�����x��a2#�D�=��`��Z���r�rbm�ƌ�tA xn�>�􅲙�YPo�/L�XB�n���@�e3��1uZ�m�p�1��j{GV�YT���X��|G>i�(>�$��L�_><�!;X����~[�B#��J�0�����A���	�A���4��/Ɍ����r���Rt���F�b��,�8�J 2�g7��2��Ɲ��@���y-	i�K��O�z�� u4��-��e:�
%���y���=����{U��53(�wJ���Q�n���'Skp��1,����O�\�	�M���'ӓ�c�L���I��CJks��4ȁ MX��?3(h�o�'y�4�"� <�# 6�IIrX��:����i;C�J�� <��O��ý2�w�-��cE8a� ��L[(i؛;�?ﭟ���{؞X4���C�oG���z��1��P,����=��ě��1A�H��o�=��Ȣ�\��φ&>{5����ѻ�<�5ǁ�<�P�Ӂ��$r��[��ey٘e��t'�k�����#���P�>���\�q�����)e�;�9|�Z��F��s�S0���P�DO����r2�� gR�>6ZDV��_�J��ͮk�����$�v��.�ܷ��1��l���~�*-�
�Js��?�_
{�
�a�	/<6֜��Ҩ���Y�}�P�v��w���5'�]Í"��8Ү;AJh�bjթ�p{Zu꽡�=���l?q���-��3�e%��s|�"ץ�-E�񸏉E8�N���0U�L2���&ɭ�/��F<��d��K�!�O05�l8��|syL��51�?���	��+��J�� �E'e�W?�D�b�����=tm��M2�L��uh�\V�w���)\B��I�T��:��VJ��B�	V `*K��z����w��?�Jͻ�nF��>l����/��G6[.��q����#�bngQ�+� ��>=��E��"MqX�R�~�7��AZ}�b;�]ްF�kw+K��J�)x+~��;����p�I�֕ȉs5���i�-��n�x㟤��[�L�t�H��Y�&F�,�ۂ���i�KA�)b�P�p�T���kK�d(0^H���,�R!�]Nw�+{Kk���+�B��3���o���d,N;�wB�5����V���=X>����A�8�=ʎ^���3B�M+i������W�f����X`q9�����~�6l� �Ӱ�%V*̈�_M�g;áX�j���^i{K���P;�d8�N�Ɨ�vb�?f�uq� ���!w@�]@�/��+�'؟	rXC}	 {̤�Ȇ�}a*�U{S��h�4�W��[��A~��GBi�+�AD�)μ�����-]�l�/l�[~O�kwQ(v_:���T`�҆���k'a��I ���rٰs+�5�4��:F�a��E����P~���5�݁1�p�s<�����'.�)�SGֺ?{�w� ��]"�%n�I��]���H����v���pg\�"&4�h^I���йr�.;q��Z;����nd1W�2^ xX�5+�M"K��Khj���N��3z�[�;���J/7r��C{�?~��� w�D/�2�F��X�6������Ұ}�r�/�D��N�����%�04@`I���[��B�+�T��#{W.^��8��v��2-�� 5e�����ȿ���>��kEqZ]�NC�ʸ��Imm��	\]#�{whƝ���?�Z��̮��y7,��w�4��K���<!�I�zT�V4>lٓ.�I6)��v���z�x;�ul�׋��Ǆ�D�P�(�SH�z<9�m�0�y�,����R0�UPb����9���&�z�����K������nK��\�M�E����!kQ_�-�fhxY��E���W�<%�!/q��eyq�����N&E�#���<�n�Ѿ@�����z#�&�^��E�[6�إ8��&�*4�\K,DɌ:��#w�kMqp�'t)L�J��*�Mx�c��/>����q�nݱA��rbʧ�jwG�E���6�! �K%�W����:J»�ݴ�x^fܳ����!u�gNl�q
S�j9��Q� }���*z�Ӂ��? ��Թ*�T޳�q�<8�:;ͺ>
,l(��A)�d���H~�)H�6T�f�]��.N-��+IҔ�Zb~J~ʌ�Ԋs!(�B�x�#�q���q��E5?B����l�#��Ұ������ң�$d���X�˵#�ϵ��Oq3�M9�J���� F�k,*a0�'8)'��R�݉/�'�ă����T�:����6��q��r�`�"�t}�	�@��2s�H�̅�od�/K�Q8�]'���/�b�J�̚���r�|X�d7�|��D!��R;{�~ރ;iy_�5p��1�@�d_�/���\?��sb}�AԵw��ۣ�Q�{�9�p�q�[:�4g�]��+$8���$���C��՟�i�*�:�*	C_�9�0��s2KyKG���&�?��A������n�Bl��8 ��`�ak�Q9���J�e�n�\t�_ιQR�6�/���E���\1ڈ��r��oԘ`9���{G����:Z'� _U�xg��WW}�D]�a)��%>�?�[�O_�\���Hsr��F�S��h�j4+	>Pwo�-��G�m.	4�_�SR��Vn�#�(9e�/@)�aY������[-��j��tJ	��40���9(��7L���ؒP�˕�(���1�OYA'�/���[aӑ�1�TrU0[�����I&ɗ���8��g>�>l��#lQ��0S�yj#���R��VWmP��˾Wg/�c`�X��4�WKX��*�^�X�^�Ȱ���:��'�_�$���9 ���;j*u՜�:�d�rE!x3_�2E�惬i_7ŭ?�r�����@7v�z^�2C`��O�_�<\�5�i>������/��؝a���
 ��5���jD^���~���ͳ K2���OE�Ư)s��렿hM��8���$��?F���3������eL�v�[�5�Y����5��a��.����%Ğ�س^��1��bW?�<�_����"ܤ'�}ݴOĔ�����΋kŊA%���WF[Y-I]�:���	9O��Ez�����灊��Dc���4�!)��Ǚ8�:�VC�W��7�G�SiK�b�.��h�w%Ҳ�-TDr7�w3Qs%x9��|^}U������OɧbR�mY#���)�I���nM?5ѣ�E��ݽ2=�XΛ���U\e�jA��YI��v�8;x�U������� gv�U���d<P�~�10 �!?cB3�N��� U��>����?;�O+Nũ���/�r��J8��i$WoX��/WV��![�w�ul��Ȍ���I)��}R�&�$2ޕ�:k+x�{����74�>�=M�T����/��.����_7���d1�Ҿ����� r7�Z���}�p�cɥ$�b�`͞~��Ԡ�Ϙ�(��jߘY�p���z�a��!<T�7d��+�f�k^��K��וN��<�3�eIOJ�f?�TZ��o�3cz%�"���iy���9c�Ip��c�}����eix������R�͔8m4��
�2��2k�
�)�+	\}@�F�oz��a���z�2�_��lr��`
�M1�u�P"p<)/[	h�
����G��,��=�?��D.�e_AĦ���VC�fU:P�rϽ����j\s��=~ZM��пtt҃���-{׽`������[\[�R������2��]����~���;k�$y�*Zi���ʲ��u���՜���=�}�d�tr�}k��<>�!������x|Q���3=�e����:��+��T'����T@��&��Vϟi[s�OS���� 
]}��q�}�&�T�tX���\)��>x������i�6^�٤ل��r;~��oόɺ�F�u�N@�%kj8��涅kP��bc��NSß�h�k���M,�l׷h�Ѵ�	ȉ�rE�����]]�ZI=!I��*�s�۝w�7��"��i}S���D{��� ]��e�K`�
��kZ rD����7;���.Q�oMw �w^.�ꕤ}����,s�o�`ކ��ڍ�z��ctB���;d�F@���ܼ�}��?e���i�q^Y����|��{L���gu`�2 ʹZ.9�J&ά��'� �%�|IhA)yp��&�|�r�����F�����Z�j�>!��q�0�>�{ɧ�h�����e�5ϒ<�p��R�r�+��8���~ay�������k*`Z����u}$�V��RZ%�;�sj��wĥ�C�<N�����ws�b[���q��3!^�xQ]�~�/�[o[)��S?�y�nt'��X�87AEK���[/3$R�7��(#���l,�q�@�;jX6+	
r�Z�P��֣�Mz�p>ȣ"�ؔ��;����@�(*���c�����c���4R�0Tp��(�]lR�P�5"R�D�iy�i�4::�=|����F�B��GvV��)�u,�Ź��8ϓ&&e��1��)B�e�	�aӶd��0�G�ʴ���}*Z���f��#Ia�M����[:@']��^=L9�Al3��LY�������x�~"R��p�t�#�ԋ��O��<��c���C/�(kuI� bf0�R�k�!�绬�Y�쭨Y��2��V5�!�Jw�)��q���9�7#\�!=NR�y���r��n�2��f�w#������ӫե��F�7�"����I>+���o��U�gT��� � nr{ 9�\��40Md�{C�&���u�h����\�+#�Dd�:�̎׎{	��V�;��эn��?�]��/�N��V��'�[:���-�B���яnK�-���1.��B���l���'�%3�uO	KC+�쓞-�rϫj�yfb�v2wt���f���Y�O��,Æ�(�[gKH��{vބ�\<l6B��$�؉6��V�{;����`�3�*���7���? ����,rz��}���X�_��.�)qq2/+�#=zʶxS1�I[�8�=-����6�Qr���Y`HX��w�dI��#'4NR30�;�^xr���Q����37Q�����V��K�$����~��Q$u��������=\�8v;s�ʈ��$���X[I�8�#|�w���;��|^�t;�0�p�9!(z��8�#��4MGlo5�y�{;�^iT=��
JTH]Mm�k�	�d�SS���3� 4e^�]�S�m��9!r}S�1/���R�0~SGV���[�N�Ҡ�C/��#sЍ*k)\K)��ʔ�����q@�J:jS`��F��]������%ۚ�yĘ��b�0<��X��ja��_��_%K�E���{h�{C�V�_ r�37�t+��`&�v��j�J�]������4��Os+�y��V�N��P,X|���^H\D,"�ޣ�=J#OCR���Q�Y�����(��z�vt|�Ux(dڲN�.�%zϬ�7�z:3kh H^�@R�_^j`Z6��
���e�������M:�V��Ӄi��RW1�ى_cV��%l��b�29:Y���K���Gb|뭍
���<��i̎�*2E�FN58�$�w_>�s5��6o:�z�<]��X_��V������:�?��{\;u
o�Pr����Y��	(ϢbA5�hwm���X��%��ˤp�٣�ɮ`�h�8C�ha<��c�ѡ��xF�Ѷ7������޶쓳���\O,�!Gei�Ǐ��J����یp��NW��<��-���Mt�/@c2?���aW��PQ�ES?����_��"х4����N��嘷ܳ;�蟱Z<�Π�X�=�s�re�vt<��q3aG�i��*ԫQgD_+}C��m���?y��x��4���_ϝ�u'[8��tk��8m%|�dԅB������X��|9d����������d ��4@�:n?YÎ[>�j0�X3�(^n�����'́Baa �z��g�/5���eH�Q��wbq�)��	��tRwl�0��u�}h�J>{&����>�&�_�O���HI=?�Zu�.���%ƚ��-^\ysرu�j�p*��7�꺍�	}O�3�����!%����>a�1y�L��&�k���@~��5�j��x���K��6�?��/��թ�2V�B�k�����_U{k#!�|�D����.��Y�h�|���저�ӈW�����X�C�b 5X��#~�Vd��%480K@`M�(��_�b��nЄ�����b=]&�c|3y���e�Mou���a��$|9: :�&/6����G"\��z�A���с|1Z剧��=��[2b��\�U����e]��`�洧`��m��¢�QR�N��8N���j�V�@yt=w���
�0�Fu�X.��sk��,Y(S�)��Č��{=5� 7mĖz2g�?��HF�_�ifop��|4C����h}��8}�	�0C�����*~ �USNy°���ᶂ2Š�jSX^��VPF�A�+�;�R��w1���^Lny�� ��=�Q��jNv�0<#�HIջL�?LT���kM5;�;��A�iڛ�� Jϕ!�;�.��=�MkM��%�~3�ڣT���Y����'�S�U��i{4)[��s���`wB���������g���VSe�������>���ϗ!`8+ǭ��k���gCnk�]r��)���>7�����o��V!E߽y����M�3���A��!�9|�\H�,�i��E����˫�2χ�k�qj!�t����Kª��(6��r�x{��1��3wY'��qs�W4��X�1^�'��2� �"������"
W�WE���د���+�%p���������:4��B�9���jA�&����vu�U�PM�J�dg�7B]��m����(ێW��q���ů�y2�A�@��F5�����D�Q�|�uK�}�����}�x��Wk��yRφ�F㔕��^()����+�!��p�&"с����d!����ʐ����T�p�Զ>d)7����)�(�H����eֿ��:GQr��	��(��jBE���H�9��=��RA.Ɩ�5\~y�i J�`�,欷fH�ύ���J�'��j���6�p�!��~�꠸�;���������+KC�s�(-/��D���yK)��p�D�:���?So��6c��.K�.�i]9���^v6��W羏oqo)�x��t��z��ᡊ���h�W瓘wR��@�Pas�~�V�en����� R[C�4z�W(˦qn�S��LZK�,H1D����� xAq-�6F	����y�{��G�6���G�%��� �0w�9�ٔ��GП9ر>ٽŬA8��E��4�Q��~w�XJ�a���uS#,J��t���Q�)���
u��)ӵ ���EKp�f��d�5Z���:��OM�+�.! �HL���,���P�5�rL�k�;�u��xxP�T������U��fp��|����6�F��v~euk�i�w��V<(�x�LR*��"�Oc����nF�����LJ5��)�� nt�.mJҁ�Y�Ze.�O*#���׽����ԍ�A*[�L텴��@h.A6ǆ(��z������"B�5)�������2JG~�뢇��fuْ#��^��Rr���7��rN� ke�ϛ%�%���IS?����8$���F@dj���v-����s_޻�����
�&�a�Ë��$��@wQ^dr7���YBe�����_��q���XG�쎠~��2Θ����P��:+8U�<|�Od�+7E��l��B�v��������	�$����tn�L�RuG�wA����ϸ|�� ܑ"M�o}�&`��!%�o�_�e㮢��J�ûK���72`��Z�1�A��&On,�K�Ej�d�x���苊�RA߷����D��m��_ߒxmy�Z���tg�M���+j1�ttz��R��t�Y
�Y^�M{��'��:��e�aMW}�� �"��J=�Ʋ��K ���N���QE��q�=���;�t����/��~:�Y�
��$�Ɔ�N�\W��l�B43�\�R��}� >�� �ÑG���/��o�\?�,�/�_92��Fj�C1���B`�[��lcY�}'D� |��$�3AB"�*��GCE/���05�-�b�V�f2�v��R��DyޒCX��c���1���,�^R�/���-xHd"I�uߺ-] ︐n>�0�5��Xq���ڄedaזs��;��=�;h=��0��, �BX=r���͹�6y2��Z�v���{R�k�-�F��7��BP����P9�,=��:
24z�c(�'D��*3ZTA
ᧂ�ZQ�`WKwY�Tױ9�+Ȫ 0��fs�|�ˇSɍ���f�u��X?�[�-y����0Dnp�I�0�Ti1jYO[���p����i��x�[�/R�sԎ�/�^�?��һf"B�IƐ�3�fhb�)5u��o"���G��	�cL��ӓ*��\�����^�wЛ7�;>������#�j����,�ɦ���PrSȉ��?YuQ�-��cL7���,���n�}\h�C����"-�� zt=Y��+B�����x�	旟f��Ul9(/?YK|���ߛ���NV��. .|+C�˵�-Ã!�'0DD�:�@w	����U��󾍴��-ƙ!)��od��x褩B�85r�/I��:>��G�bMգ=���̳��j��K^�34(�)���X�K�W����rk�����㫤�R� 7\��6�Wo�9v{��ٶ�q��²�H��u>v���g������#�b/d�}H���!�B���U*��>OvM^�j�sl������r���z�E�.x�9T0o�6+����d�Yv%]]!Y�����I�h
���\ܺE�.o���&�v-�d�?m���d��F�>���u����Qס�@m�#㐐z�*�Ɖ�
O� O�e*�w��tW����S�8У�dpYz�k;��a�
��26�]��=u������r�[�,a�2���f{���f3c�Lmf2�pSr/_ہ�	R$b�5�,�v=�}n'�wFV�:�a������ @-M��;ڽS1��p����q_�޷l��[ w*�@RC�`������5'M(���������v��kT�-N*�j�҉��p행�x���7���o�>l���2H .��6���d�kRSX�K{T�F8�_�1�TH���QD��$�,�'��Z�i����#�2�p�b���i8{G]��W����+�a3�?�:����i�O�	\���b�Ϣ�\�T�ڼe}6 ����A�'i�	�^Z-,CQ/+$� j�Q(���sP�:e�G�ܡ��e2Ța0������j���f�%?�/{t̀�9\���<��TX2M�f��K�~�~�� �v1�����n�H��"�e��Z؎��l�s�ꂓ�!��B~�)�srXEf���$J�E5	3�q�&�?�W��{*��%\N���	3���9=�WN>=�cQ�c?Mẗ́��}v���6*�ea������`��$ ��iC�G/�դ���`B��e�07���*:Q�r;�����GBݦ:ʎ}(���  ��(� �d[G]�c�O��g{a�5�sg����l���>�(ca��Z�S<�1�L+G��đ�z=�P�4�)_�[t\��8[z��Ğͬ�>_L�o�F�����}������Բ[�2����{�٬�ڰ�'����GpA���q[(����M؂u��a�L ͅ�t��/�R������)N����Bc��b��f��9��l��'�[��U��X->I3���#O��,���!{;]�N��	d���~O6� ����J<}b�Y#X�g�GBa�/@�$j0�r�	Ȍ��*!�ز���]�����,�t.$o)�p����>��RGv�o�yz89���XH�7��q@CMp���F��
|r�����h�ԉ"S�P G���1��-=<�W��
�!�O� {�):q����J3fF�=�Z���w���)ka�BSǱi��y��f���Z���~�ڌ�0tO��ێ����
�@7��e򪩴�B�p�Ƒ�;Џ!3��99G��}�kU���UO*}�v��>����F	5;~�pü��(�ȟ�m�ǐ�?�IEL�� �3�����0�]�6���qCQGG�y�&�*��*�U6���	� �}��	��a���:K���x�~0|c�l�qx�G�z���g0��`8�&����+<��_>����)0c��/�!��.�J��[�-ٚ$7uE��Y�o*)eS�};R�����/�YY*lW��=Rja0�d��!�O0�#�)�2�C��}"�̮v##	�����놃lWBx�z^u�4�n��@H�F�q>�Fc�CP�'s�lᑑ)�%߿	����˰;%��yIւ�EdA��dZi;�楰��Z�njb��{~kd�	�����yY����Ń�����L��dL+�x�H�(s�Ѽ��kO"S��0�$ ��� ?HE��p3�I*Y�q[���Iޢ}X����2��M?a�]��e�UF�M�P�'G�x�����]��R�����T9���&茐�E�7��פdr�w�E�֫��_Q���v��^��]�a�<f��lD6bH��Qu��s�-G�$�Eэ4�l���Fyֵ����C��s�}�q��]��鞹;
�2�T����I)Vا+��eQ�*]���FRB��z���z�%���0sT���saG��H�9���Z;\GIB�.R�e���{O4�2�!6TwR����M�˱��J�˵�k�1��l8,�k����X�:q���r�9�#�q�4O���h�7���L��'��ި��U_ƃ��*>rL�ID7������/��e�re
����]Y�r�oQ�?vm�^���M�啌��l?���~�h) c'��(I�I��r-o�|�}�3\vj�����
=]�9Gn�|qH�MnB��_ts�`Q���4]���3���j��h�F��3� �}�;,�_�ByB|���|�[����y�Z�~u���)��*2�i�`�Q�XDZuB�U��xT�2&�ρo�m�j���R���>pA)&owջf�-��N����kI°^W'Ƽ�E�%�-����*���!�����XM���b�TdF����tۧ>����;��i����P^��ܝ��A；�[�w�rN�ʶ|��.Sb���c�o�V�_�$�咹�?}9��8!��[��q��J����ڻ>���r�a���iǵ�s��!;DM�$���{�};++M�#��\*�ݩ5^^�U�׹4u9�"2,���{�R<{a���-�V�=�/�~/�����ރ&f�� ��1�1�[n19��̎	��d���T&�jKw6
��9�?�,+~��D��z��$�� �{��a���c�wPOc��B7$�gV������l�M�j2f���TUv�9p������c���6e��!��=���o��m����^�Ĕ��x�{%���>s~Ąa�E�2c���p��qջ^������ߐŀ.�� �c�j5�qq��r�AAri�-���^�4��i��R�%�G�M�_�;ϒX�c��@y�6����4�.���0�ɔ=��Ռ&??�����o���ō}�MJ����	����C�ZDL��������C�^�b�ؓ��>��V|R�˝!6��?���w��Ȳ���|\���
�²n4�?1�?�E��d��������l��.�`����zL1x{[�+,ɭb�-���X��0��!$�p�u�'�AL�."(��L��K�k���׀�l�q׫�pj�>K�xI��R�S��e;�A��3$�l� ��V�M����5tҠ4G�%bs\6�<6�0���[@$�:̻���D�5{_�	�ȻI� o*p]yy3Eԝ��B���E��y~{Ћ��9�_W��`�Kr��J�.�*���H�����_���w�p��a�/�C )��Y�Ơ̞�ȡ�r�i�E)t�Bș�x�ڲ�Ҍ�@W��\|�����+�a��H�= ����<(WQl�ls��-�HI�W88)���{���An��I�EݙV�k�Tw����SNr��OP�Q��C� k	D�v��a�mO��'��AН��2��{�d(g�����0#����U�r��/����';�5�<�>��]vC$>�Th�6�*[
��x������ļDI>���Yp>�8�B��6�n��jw��qgs3+�5b孚�?7r��>�=����R��-�`���/7+�E9:��z�ٸ^)�^jd�j��<�6��&(���+8�qL��1�@j�YD���%u�S�t��&��vA�(��0	��u����'���7��ܮ��CF���XYN+�N�f}I|����W��I�8u�~��Wq��_e658���c�Q\ZB��If�F�۝/7�R]?�1@��֛*f7S��kc]�Sȸ���4q\(�6]/��I p�Js�F9�X�ͽf~6�\����	@V�����Q��܀4�|�1��&��Ҧ�U��`�6�
�Nːl%�K;�{z�Q6�vċ��_z�P=�D��S�{S����l���B�7������f~_���M�b�<'��2}�9�i�Qʀ�P�LH�����Y�)�X&����S�Ď���L+��E�L���#���X́�ULmလ:�@��񺂷��Me���ܾM*̓���6�$]�7����a
���E2���P��s}��[l�-JY6r'yRk{[;4�����yɤ�F�nDj��+�?XL�	�욚/�li���i��ѓ��{۱|���0����N��Id�|��ͲO����{V�N��).�H�\�
EY�^`M,�x4`�q�� >��Ʒ��I�^��?�E�n�7� Zu%���=Oag�mV�Zpp����q���/�Pz���3P)F��mѻ���#�����?�����VN��-|^���}��n���Tb�W}���t� �B��,ͫeFر�D7�mKm^*$=U���P	�|�u*��Q�]��M�v8��s~�>���J9�|��lUV����Iٽl���WU�Hܛnk���#S_ewNs$"��Ӛ<̭ >�E��o%\dX6��r�Q�w�"��G��Z������_D'�;1�~����]E��qU�d\}���Qd�_㺐,��{$6�+P:�M�E_Ӝ,�ad��>]�b���]P����i���aڼJ�m�0� n����y�A�hׅ�i*�{���lJ3�&XƝ��U%���J{����>~ �n���?��+c$��_5$������0[����K�W�A�\�Y3y��^�_%Ǫ/2��B�h�����+��C4�.{:���1�j��g( W�~�{`� .&9�խJ�C��݀Wu\���4�v͟�g���,Y�{`|��(���M0@Dm}^�B�(s�Im��8����s2�ӄ�a�mU��#��;b~tz��/ը�[y�α�H{M�+s#���k?��Mnss�P4�Z,�$��cu�l����y^^怯Ώ����u9
ą⇝��]�~^�g��?�,`Ai͈�%X�'}�*{����4��:<ҕ/M-����B��\A���#hj�@�R���NY.�l�pBSN�Q�("�ރ��_��W�y!��v�6�|#X�T���QS���w��XaL_J{�3��!��р/ʏ�˵зu�h��w�z�,$���)�M��{O<�EN�K�Ҹ�l�nwއ�n�k�ܞ��G!�F�gA���3x� t {	Za�=
&9,�0�����Yk[��������H��R�?[���-�H�������@f��R�;��{�f&���?�7����ة^)T��-)P޿G�u��m���n�@��Y��Ň�����[J���K����0-8��D�0��LlH�l䧘�é3y���8`<^���f�)Ϭ���N�c���\�R��f�l�X��b�e�jYT� C�����TA�_H�UV�؏t�����r)�4�Z��	�9+��y�K#�7胩s��r)�*�t��X5�N0����b���d4?����z�B�i��Pغ��^�W�����'_�D�M?�=�
K�["�WT�$�'˭ʹ*�8,hW�G�]6}��>rw����n"=:�	�P+�o����,آ�/��e�_�G-��O0GZ>Ma�z�mi�V'a,�I�,���@����b�Y�~Q��8�)�@��c, �U.Qy}��<~��oz����F�)b����w��X�uQռ�N��\$�0(�v1iҔ��V�%5�� ̋j���� Ԃ�V�W�*:��~N���X`��4g����w4E����gƲ��IvVXYoT���Ed�j[��n�4P�L�_�d�0L98��@`[O��8�<�:�l �]Bܴ�|�3�N�Vi��Kظ�Y�SIlģ�'+J$N����G$~�K\��:B�:�qȝ�S����
\� �|�;�q^+����/!�j<�\/�7d�T&$�����9�ì^ꮊ����������7�O�5�0��+i�~kv���M`ꍕ�W��緉Hݠǵ�Gi�`��:l�&�p}�%���:�Ӑbũ#&���P�e&�a�����0P×A�$�c�y
q��Mj��jy0E���眭�t�.3�H�"�4�+��a�\KdB�K�k�pS��L(��i4�n�˙I%�CP� ��R��2/f���\y@�&�׷�tx2۹�K���fw#��6��p�@�2cJQ^CGŏ$ �|�U��MhR���D:/��.��F\Dr�P��v�E덑��NM��8����!��[0���x$�	�"�q66���3n5�A���.�]�9�S˕%���W����.�$�\��U���`�! �ˣ��r8�G��wz=���m�Y�?D�p��y������N���I%���6�k�Qs��&Qz���0=�)y�3B�������
R�\7T��a����#�x�ba�-��s,f�;�a�ᚄɲ?z����3����Ko��lCO�؎��Y���J��El�ut����%�]�I��Wq��� �ا*p�Gp�Ӕ3��|��'���}tK����(}�x�4w/G� zg���!d��\�͜��YKĨ�&󢣀j]^�w�<V��ܴ�!^�� E�Ƿgd��c��w��tg9'�����K=*�CΔ<��y��������ԢQ���*���B(�BEZ�%2������h"7\H�Z>�!�Fc�m�O�F�硦�2,�~)I|,dؼܿ3�	�D��=l����)�Ƒ��h���c�[W�%��(��M��}|B���'0��B�z��L�O�
���g�c;2lv5��Qn�Ɇ~R�IS==�Z��o4G?DpE.i���he�c<Ԙ�J}�N��6=�'�Gb��<As�0 ���~}���1a��f�@��ʕ��ގ�����Q�㦤'�w���ҵ�Ls7u���z�g_���������h���35�����O*�1���l���"������{:|e����׽e�&j�2|ꚇ
�˿q��R�/ok�o�@�f�X����W��s��q�,)�7m�I�p��H��|'��Iל��s��x��/BQ�yI�n:|��(�]=���b!R���R/�2L��ެX��Y:�6,v���1_��6�|_��;�� "�䂁�#3`���)sdb�
���7�y�4l�㳍�Oes�!j�(N�̍I��[�v�K#O���w�T���q~B�( kY�� �[����͖���=v>���ǈϲǼ��vD~o&��|%L6��DVŪ�Y�F�����WМ�k �WEJ�����O� u�Jr����pym5�F'1p���"�g泳D���T��$�<�/
D�SQe�@�YH�A�O�N���F����ߵJ�Ud��J��1���^@�3W�Dn[	����o:1-þjv��{�A%��жG� G���:ye	���kwy<e���C�U�L=�9y�h��L�d�NHO��&��y�M`���J�[5�=h�|�C�zO���x�S&�J07� �fI�6�����PJ�F�E�-:�'��4l�xtU�P�}�0w�IJB��m顩�O ��c�#�� -��|��;��4_���E2D�~�oI�U���S횵�*c-B�d|���p*�=��/��LB�߭�k餩�h	�ܤ}�%�����	�q�W�q�f�s��A+i�FE�y��$��ꨝR�������0��z�H�̥/q��z��}��3 �l�/Y��"�r�ն0o��~���f&��v0��I�T�� �'�m�����Ԥ�7��^u�pTOǥ��}\�)�g���'��[�q��$&೎��D{wT~\�%�z �1��I�h��3�R���8��Pq]�>z���P����Fm폨��Yy�����Y����T��f���3R$�t�NkgMn�܀_`≑��!-���EO��:�{�\s����NG�k�����QTv��z��`!�{�,�� 熑��`��q.UOy-�,�O�4�C�]�5d��&s ��\K��M�!r��f�μ������3*�
�4ebzpt
 �pǢ�F�2X�v��z�$��$"z�ۣfl��!�Á�&R5���Ch����FB�D��0$ϡ�U��ܗ���w�3P\��-Nⲣ�6�#r�cY�
���v��y���"��gN+^�H�fӺ�$�uΉ���x4 b�]�)����D\h�Q	�t���c�����n�C7��������1a2k�o�h)C�p��9W[r��6xE�����_Ci��λ�?����670E4K���#��g-�N�h���s�k���� 77�+L�uFNԖ����,[��~����NX� ?������_��ս[�hO��4Ϲ�t�G�~�[�8��!ȯ,52�ŧ�;�&���оmٷ��z��-�K�b�0�ۄ����� �Cf�_�:�>�J��H��	��fI�d��\j�t'̉P��NO`�'��䢷R%!L��"����AB1�JhU�'ۢy:X+�W}���vD4A��ثV.�go���n�`P�(�ξ��  Z�H�$�A>�~�ۋ�[���}A(C����xCp����گ������.D�/��#L7ϷV�i��|�*������ٺ�����sV���Dr-�K��r��h��E�k�+@b��GH5�m�ϒ�(��/��I�F��l�nV까}���qwIK���7=�č��+q���Orz�26���p�z�f\���Mo�dC6=��c��֫9��)����"3��m�7�Q��@�*4���a��V֏pǢ�r��v�c���J��L���{�}���E���|oob�M�C���o��a6�h�d��r��߭F�7���+�"����ر��ct� �e���!�P�6�a�ͱ�[�3:�
'��ԕ}�)z2�rc��q��΄pX;�4�+�	sXe�3e*��6�+� V�k���gd޵�g]�s��h+emԅ��n�r�_������=��,� �;�j�����n���퇣1|�:���_&B��j�v8��|�M�K!��M���e�=U��dA'w#T�g���U)�dA�ƅ�c͗P�>PHH����(si�c��!�Hձ��n�B��ߐ�}����x���مcf���(DQ��%�ȟ�GW�����V ;,rG�xP�4R���R���ooT
�d�ݢ�0��SᰓF�D�^���-r���w@M��m�j�v�M`$ 3�
*�dE�W��^|�m���W�����ڑ���(B�}�>�k�9��x��/����Wn>=R%�"&���'�Sn~v�Ǉۭ��e�!4�� ³a �kT�;�W��ΏR�\���R�o�@Y�tl�+BΆF�xJ�ɜ�	��M��$��Xv�z�$�fP
?&����TWX��B�Z���~n~jO�1s�HЇ�S`�#7�W�dv� ᫌ�ea�o��KVP>e|i�!�dws
�hBL���Z�i1��:�y��6S�cu1]����F�a0��P����#���*�r�l��Yz�%=��71B`-�10^��)���V�r�M������(�
V\�er-���6$�~-��3�T�����&0��^�>��@y/Z�))��UN���nx�$b|���Q��o+�O1�����M���f�c�^%vߒ`��ȳb@f�����6J�~ߺ-��$���Ⱦ��1 �ib7A{��)��-	5?�,{.��.���׭WL�Gx�8��?����[,����u�
�b�܎�hګY'���ϒ_��#��C҉����,��1/�
�BdG@�;�?Y^�UF�Ocp�Z9(��Ĳ��&�͸�����P��sd��8�L@@�������H���B�(�G�`����	LAЛH���BvZF5��� 	�)0��.A�|{%�����Q�DDG���S�څwJBp���s�A/#�7\���L�U���|���%������=�P�Q�mR��i��;��˿�bd���{�����O�$�ɳ#c�f����h�K#�.�yV7�R��e�H3�ז=^ � ӡ���b+�5_,�	q���Ƹ��_cnE���ë�b�!0,�����Υ2�����r=�3�����\D��G�	�k�j���p�q��-"�3�Me�M;�ʅ�8F�
�g<Mu����N��&��pN!�Ikt.#��8��1k� �2\����$�b��U��^vo6��Č�1�t�Z'�K�[&���������s�J���������T��kǖh����fi:��e
�8�7�O��]��+ S;'j����7��i���ϭpՈ⬕R��x�H@FB'���+�۰��t��9`�
�UJY=A���2�p�2��1��Ҳ~�R����n.@�Q��"d{J0	��Ik�\���4N<��~w9>��?����غ�8��80eմ�'��>��>n�����S��lh-T�lH?�S�xG� 5Q[5LԠ��db}� ��e���=F��)PwG?4�x��z���4:�p�|��|I���D�p���N�6�Aa�	wӻ;RP񎤤����ЎH�6�Ѿ���f������'��o�0A^�IyR��\�}�O=6���ߺX_>�;.|�
�u �.�KW��o�E�0�q�ܾ��܋���X���zFy�~U�.�x:0�)�� Ͽ������左�N<a��I���&���@�~='���X邊�@�5{%�
���Ő��5�@�(K�DC�]�y����0�f�N��	|l ��۹B�߲��׫iL�	0��f�T;�T'G(��Ɛ�}Ι7�����/o�
�}&��"���#9�"�hU�d j��b�j�WE��L�9��wć��4d[��jy�S�p?sa�VL��Ͽ � rяhտj��v���I�����\Q�I5��t�� o�%�ɒ�-�׽-I[����0D(E��'�s~<ෘ�Ĺ��.��[Ru� �v�kP���08h��Z�63�	�^��*B`�i��؄���������A8�x$Y�5v"���H^S K/�9��ZŉP��E�f�4�x_=��ȼ�{���5�RB:�9��B��Ы��󃳼i(�Wqg
%�y�l_O�$c+U��ȬT�.������y�b 뢎��J�ùa<��� �;�iW֌Q-Uw6'B����F�q�#T���)liy�y��:G0ݽWX��[,��a�ݏ[]+��줆��3B��Q��u��/�����%��w�C�˼Si�	�&�n-¨�#�O�G�쿊��UнL;��"�|<T���4��Ǆ"EW�3Jr��K��/:,O�k{�i���wRd��.��f����Ws�e7Mz����U�7�O�f�*c4�T#�RvQO�g�aLH_��'�#>�����T'Y��aF M�`�@O��-�p�dTΏ'@]�>��{��A2�@"��Tg�1K�?.���Ī����Ͱ�˯��Ȉ�L̃�����2nd�cե���5�7K>Y�Z"`��G��p90G*P�Bf�r�Y���XaKМ�ؒ�p���
�V4��Ռ��U(����V��>_�;-yA!��JY8ve7��F??Y��(�����|��qoAO3��m\�tM�[��!�i`rt�(_�?���!�6?�s�Z�ʟ�=$�"i$��]N�71�ټ$�4���3��w;R�5��I�� &�Pa�C\ws>d�	v�>q������A$8/a��U��9���/:7+�{���x�.�����}b�kg�EDN��W���K�^O����q،S� ��ž#�Yt�V2	r��M���:�;��Ie�Y���HR$�D��b�iR��RV�(���<��,r�a��K6��u���0B����z�t��Dx������*#�ދ�Ovc� �������������%"c�Z�_�V���V<��։�B]D;nK�x:UW=@r���o�UI���O�z@���0ub�c>�7�>��i�lP1X�'�9��`��������ueϴ�;%g���<r�ǡ=��<i�Y�cv<�g�)"MfN\��R�cU�MvJB�
)�u���'dM>�@�,y��Dg��	� �w�:;���9���8�1�=�&�z�w�2����{@�ڛ�?3�A��~W>"�����>�*ެ�I����(���8 ���,>�2#r�g��\䛨�Y�p��۷@�X��&��4�L��}�d�O{�=%�?�hn�N&�H2�w?&�|�L�q����܂�p��%>�'�������x��M��sz>i|b�I��4l*	h������v�"���P6Q[�[Q��c>��mh]�}�햚�_�ۊ`��^g��ฝ�k��w��.K��o�$U�7�W��婮�&!�>������������	�R	Q��z�7��',���.-����Շ]i��R�%Q7h�A������w��̥��(�ٵ����D�xx�/D�����H��iR�k�oT��?\R��m%!,��&1����LU	�?����q���'ϖ���ި�i��Ƥz��G�<�h�e�aȅ������_�9*MQ���>l��N�H����;�I��/f0直\>>�J7����+�@�t2f#2�����v'�c�0�<��Q�*Y�n�~Ҩ:��ǫ��s�L�h1���G�3���'%QL��E����K�$\��i;ˡ�f9�u$�{�b��K:��ы����R ��R�{֣Bl=��+2%���� �f]1�4�H��g����e�b����AdWT�O�yȫ)G����{���0z�Q�]3����Bp�>��#,����̸{�K���!�]̏@��Mk�5/����=h��'`ې4�������$jԊ�X�a-�	ei���)�uY�m�j���hI�r�~�_��n}C5��ؖ�E������3�c�b�y~�b�L�r��֍� �N�$�N�(>A`�jmwx%I$��"���nH9!�	E�.�O�"�����3��g�_$��`���{���u;f�!��̮T�����{"�6z��o�%�	��|�8-L����	�>�/����`ޫΧ�d�0\8y�$0-4ݶ9qŊ2���Jx��#1i�f�t?1)Cl?P�4�	�����Ji�@���.����
�*�1�`u�1�L�<C�N��s ���鲿9,<k��:�^�P�7H��ƚ�X&H(��C��m7A�V�N��'[�����H���h����
?f��ш�vB#�x\�ߖA]�f�QL㝳MR�s�T� \��ZޫG�" �r�	�����+f�X�ĉ�͈-h��^Sռ����w�ڝ�&��cÝ%�;����J�$��w|ɭ�Ϣ�r�s���R�F�F7��	Y;���9
/R2�M}q�+"������� 7�/}2����B��x�C0;=����VϮ
�_�,H�{��x�>��V)�����'Fh�R��������H�����m���Sj��s�&?n�D8*�-��}!��3z���S�,�f�ɡ>�k��*;<�����V5�^�#71��~�yy��?�^�r��YB�<���{���xu����;���PS��X�0h����kLm��#��bx�=QHe�Ƌ8�������B|��o�2�ˣ�ԉ�Ȁl4d�R��;�eٴ�:��lj���'�T�okӊ�"���ݸ}.� �c�k��.� ϙ�1,�O��G*ZԹ^)迊�7�4��"�z�^�b۫��d�	�i�ո���IL}��H=��	���eL��\���'��0'@g��A͒�b)��|XJ�7B�0Җ����	�����d\Q���V�-?��ý����K�׏�&y�4���y\�J$���1���=$�b��<
��o�J@�@�O;���z���8_b��p�8�Tt���j�) �KG"X����ޏM?I���-��Sb�a�7����Eեq'���_c�xvMƐ�xi�?L�±���X:Rb�	}����wۚ������&x-JC���#h��]N��-!T�c��\@(l���`�Sĸ��ł�L����2�!�h�:�=!�8ג�I��`!����@�P9<~��c��Ʀgo����Q�V��|�N�zM�S����a�V��]�1��w;┬�h�B%
�sJ;�E\ϕ�Ϲ�����M��A�&�m�:>���䲿��4s~L�z�����B�E�5w9z�;��Y0l��E����+���馂@����H�e�y}\�
S)��u�4�W|��VF�Ts��³�0��9��ȳ��.1�+\��=��++P��������29:��`���-����q���%�]$�p>��|j�0��~I8f�}��m��(��Vy�S����0�YiAˊ5ɂ�'S�cɤ6��B-���0��O	h�&H�˹�wt������A��ԁ�B�s����� �=�g��ϡ9f�MЭ*m��%L�8k��e\�{@����/F�nW��t����Dдz���
m��D)�ld�N$V-��4- ۘ��
��)���Q�?�����_1�,�w~��i��9id�X`��ϻݧt������[��c���2M�EB�5�H�Z� �Z�w<��Pc�P�$;�@&�ȶ)�x	g��6� �q��ok$�Q�4^(Ыw�-��Z��(%���`X�S���`��a@� ��a�xAV�"p	��XlO-�Ԅ�����b:�l����,��?0�r��� �<�)�\Ӏ���ԅ���xn����}�*gHko�[:�ޡ"{�%=������S7���t5�V���{a�J�a�S�q���E�y�ɫ�B�Z���mt�������U:O<��Tt�G�V�t�� �Z0d)��bv+h~d���>���Vx3�(#v��q��,��{��R��M��3ԕ�5:;o�O� �E�m�.֥�q\�l�3V���c{a����\��K��1�K�
�Z�}3;���#����cQvU����~�Ի�9+������9ɎU׻q�V4��ѫ ��]���O���(�.6���e�����{�S*i�3�ٟ��z%����w��I�1]i��*W<j����|sȁt�#�(s�WTH�2n1$�"���)*� ;���a0�î����X
�oF�"�/�S�5]�h�p�PE�P}��:��h�2��3����JK�Mc;�b6�Gc��N�	u��A��G'·����m"��,�PD��m��`��5���e�Q��cܷ�䃩�(�M��2�l�nuFE|�gf<ٺ���+�T��X'q�}	�!p���<�^_�$�jV�3��ƃdى�jq�W8��YKm:�hXB́�v���K}�14g��[���N�3Z-(��>���&L��r9U|�FH�\C��՚�L�{�!<ښ�Ϗ�h��]�YR��d�Q7�����܉��}Wy`a�<ˁW�S����a)f����7�A˥T5P��FP�Ϫ�r~0y�/[��c]�?�n�Ee��qq��1�&�����V���<�ꌪ�j����O����OZ��L,�L��� Kr�65a�%��e'ˢ�eZ��{�*z�Hm�z�p۪{)}���9^���2t�<��4�G�Ԩ?�xҾ)������^S��KѡJ�*0���#��7�Uߪ�~Ϲ�*���sX�D�����#�lwa�"� ^���^7Z�
$����u��e������3'�%�<�b �<�*;���n3ߧ4�K�Dm{�O6P!�d�R%O*���"�*>C�����{CS����Z���c�*�\x���� �%4��"k[���D�
:X�W��?�����c#�r�?����CF�'����-0Ƚ�Ü�����oFȤ78ݶpY�/w����V��(f�y�A3����".r#\'�?�k��ъ��v� �(Xb��0dI0A�"�����s�k�PLWA:xa)��Y"�-�����o=Qc�Q���<�F��O��l��$�*��?�J�)ޕv�N��6���ܼ*�AƊ_\�H�V,�m"}�&89���߻��T����:�ݲ˴�zl����h=�)�燅�o�Jc�M������Y�v�o��"⵺��Y��������9���!3a14�?=��=	+.6�I�_����Gq��UY)���+N~VB2��:#�04i/�
�AM��T>��~�� ϫ�����@�H�[�X�&QZ������ޓ��ClC����ؘ�+�b��q�a����7�l�H�Za��Y���Q��F?�Җ����c[h��{,M}�H�j��^���Ϛ��'���2��ף�#G���烵����(^����ԯS���
E+���Hv)���t����+$#ES�WM+Q��Ӧ7� c�a]�a�)�z�z�ڻ��Q�Ȼ̣�'�bP�.�����6�i��;Pz�ڟ#�w� �"�<�����N.Ő����q�?v���Q�|��Z��&�`��O�0Nf[�5��x;Kiy��;��ƕr32z΂h�w�� ��`�|&�-��A��$$X��,!��Ͻ�{X�� 2��H���q���h[��^x�g�Hy��l#UԶ�	�u��K���V��;����;�4���K^nߓ�[�Ci9f�Nݫ��Ywxy��0���B)M�>���>bq��$Q�)��y���Y��ȹ�H�˺~ghs�Y[� ~��5a���޾f9)��M�lm�����SY�Mt�6�$گ��n�p����<���@��G�L	֍�i��?h �8ub����t'	~�H�1i�J
H(��[r����߃vG½�b��VkQ��/�R�k��]�>8�50�e-���8�iB �|YH��ll|8zB0B]��\匵�S,`�0"A����:�Eh��@��v�G�ľ�?X:+�_����/
��[t��BъS#��A<9I��m�+�&������B��^����6,��5��Ek���6wvfNH�zI���v�,$���ڐ�(2�s2�_��1
̆�a�l�x�#�<e�����}S����P��eٶ2jT]��H�y�6�R9���v���=E�<���0@́�Ǎ���a�� �IDy}h_y�͓��Ip��&7��-�8��xB�lz?ε���$^!���G1B㼬�5ɬ����b��6�Q��O)X��/�q��to���sԶ�/��𺿻�M]�K�D$�N͹37������23��Ȉ��i�N���׆�����tF�X\��''��F�=A�Y�S�F���rz631�f�f��2�6�aI �Q�)p�$�D�ǳ��X��9fXj�e�y�sJ�Kx��Ā��=^��8Z P1�����Is�W������aN'3���BՔm�{B�7�WdN�R������mmz�������ݺ�ǡ$�o�>Է����n��g��;|�>��'��w���U`�z��T���Wzl[W����N��M��m��ړӈZ�C;����P� m<���K��i��OD!�'G� 'Vϐ���� ��z�	H�1﫧�wN�҆+���ϧ��X�[@���	�ω�юM��[��D����������޶V�w��y�=��)�b�%o&�#.�a�r�ċj����FV�[lp��W9��5���UW�M+פӪx���665�[�E�^ۦ_��V~��%��ĿR
h%VAIH�ތW?c2��p"�.����Hr_'���f�8(��Bs5b���d���ہ&�0����zO��^}��_R�yX��|4Rzo��qN�Dk~*{���#������y�� \ڿ^������{�*���.e�)��D:^*�u�KG{;3��Z��V�eȓ "�I���,[H�bI��� ������4P����XǷl�I;塷i��r�R�����Ri���������ID�1y�t�I���X��W�'��YAx�`��FA~Еy�^^��Q.���Z$����Ω�yCe<3"/�GU�cL|	j!���t��F���hJ���jB������(y�7Юk�,< l)�I 2���n�i��[.'�[$Që��v3M�'/ۃh���?ɔ��
wı^�niq���>���:�.Sе�t^��E>f}��F|��:1d]4����yH��c�����K���(�o�%kZ-㞶�m�k%���cuCD��>��]�<S2�f`�=3?�n�lXdJ�<*�q{��v1�xm�%+E˫H��A���$!J���1z_�X
�c:p9s�K���V��X�vԱ�������l��	8m�Ń�k&�g�8F��7�������O� M�c]�+y~#gX���`�d�t!�t~�#��c��&����dj�������lG�	����bz�\% ZI����mh�f�w(�y���i4&�+��/�$=7y��ǫ��o���q��x�qjľ�i�� 'y
�,{�+q*��j͛���E��X�IO"��L"�-(��IT��Ǥ9��L�ywg���.arq������ēs�u���g(qT��(q�4�������J>A�^,B���9�("���92�JP���چ�.�"%�^�&*[	4�کD���<Y����]��_.q��6��`ۦ���W��Hl��O;#�/�qE��_A)?k����K2� �!���s}Xn~�{h�6�:�˼��l~	?��7K�8M�Nu ��\"����SĪoJ�S�6� dSŲ);R�8m��G��«g�u�o�AIE��ԣo���ك�P��=�����0�uI�T�!ckQj���b��a�8h�eÆ_`��e�Pw��8ݠ��.V�ԫ����%"�MQ�=F�N���Z�����U�~��|cS�v{���p�;����b�a�U6[�U�U���U��{zw8W�5�PB�b�=x(eu���F��e��4�8I �`4���Z͙�!�n�I Dw�n 6�Ap�����W����?AnU�Vs�Ʋn���A1��ᶇj��7�j��(/I��CY�&C�b޼ĺ]�+F�N���&��G>��Nؚۡ<jM#a��m4��@ � Y/��CP8���i�.l|�V�:���m���|�C������m�0����,��g����4RJ�~,<�������#�aW�
���z���y�R����aUZ�gK�|�g����>��х��6�G����K`C�2�Q=f��tz�G�g��P��q[��/��$G[�,��,G����;|�b�{�{|�cՋ-�;�x�b��Y�{m�ψg7퍚��V)���=����w��P-�	@7u�X��؛n������U�!���Td��w�s|�IqH��ʝ�lwRT0:��a��+y�w��a0-ô���k
�Z����(���s~�o{c�W�eU�lJ��V�<��dJg�|SԽR[|z�t�?�	ƭ�s�gSC<'�Bo�ie�`6�~��Z^IXFofFn���amb"�p���)kb��+�v;�=のK1�u`W�����ި�o �X��O"���;`��i_��a�9�,o��S�%���L՞�R�s�U_"�;B%C&��"�5t���`l����V���9�S+�'��^p9�6�=Ri�(ݔ$�xH��ST�>v���aA�ı�*�I�3�iu����>^p՚��G������o%�����ۋD��<���>�#�T�}4G����U[ȓ����~_XG���n�>Tqۿ���m��gA-�#'���p�Y�ﱩE�:#:�ZD�S���pxS@j�B����~ȣ��'�!K�n}�,�����g�	a�lI=S^aC�b��?]٭|�A,�Pdf�ֲ@%�# �;� �srݗ���ڠ�nΚr�E�[��@�ɘ;�洐yPl"�-���y<D��ﴀuX�p$V���4�l�����'�b�}�`�&�6�(�hj�D��_��Ah{+I��d�i���/�I�"yA@3����j�qѪh%�w<�L�"��X��j>kU*��$攫��*��xN�u�'/��3�e�IW�%��e1���똜B�j펥2��IJ_ڠ�� ��r�!�^��Ïm�Oa��[�8o���Q���R�@x�T��	U���c�];gY��o@On��[�LC��k��W �X䩏��|0��I����䯨X�|��1�`����ڎ/�R��X"^_��Ւ"ԗ�{�KcH˄���| �y�D`��9�a:����۝c��;ʄ�&�ZH.]F�?� ��k�S|�}�;e�2JU�?�q7��7�+˯o+	\�F�N�'#/��ܨ Cj�.؜}Yb��G��ه���pѽ�	.6�)'� k[Y8��0u������QN_JD�8��@�uґ������NP���VH=�xf%��^;�/<�$�*���{9��G*�z���H�+p�����]2[�R�^��6�;��tA�'�;�i�\}�s��29{��_�KLz&��P��j�(=��T��)��`���iFJ�$;q��_�h~�|�ʐȗ�]s6yjCtwS���@!�m;���7�j���j�<w��nIZ�s�ǃ���ֵ��� T6���[��#Be�\�1�ȹH ����ԏ���@>EzK�N{���M��8|!�Ë��lB�@�-;�Z��J�M����������������qX�%eo�@���膊�~{�$y�y�^0�-\���I:j�l���b�k�$7��Ɣ�5�oa��b��0�H�L)�5峨�b3NZ���OC���F  �S+^�:�7T��{����1�f~�L*$��ƥ��%ƻ�H�ȷ�&!�,�r'\/*)1,|�N$�+i56�DZI��m��Nw�7hH��Q�(:�w��hr����*�r�L�Q�l�����$&E��A<Z�S#*L��أ�5y)q���ǀSD�<�8YI�S�+u(�E&dSιc �n��T%��L�j�?�k�2C�~��k�3Ms���.Ȋ|v����ٔ�AK5n=�hQA}�2?A�rU��[��Dϝ�xhc ãu&����@_�E���}(�pn
�)��I �������U��/W��?�E�K��L*����$�<{4�#t<�X"�^8Q��]w���j>��Q��R>�w�Ð%�r<M�L���b�WW���� s/�tC#oL��/였�uP��,Hj*��
1Y*�F��3'ѧ�����?F"�1Y�/YOW�)�'rl��N�2/�t������L�AI�Õp�K�X"��kX���B-�@=qN�xI9�bö��Չ^nu�;۲��b@]�����������O+B�+4��x�61v_�[�v��}���f����$b���?j�hcKU^u�'Ʉt:v�1(�".��>::*�N��{���m�MMȺ���y������<����O^kB'9�l���~�pXɅ����[�A�8_���)�I.Y-BW�X�
JƪH�?.q3��X�D�$��]�)]8��&X�����k��Z��7�`���CG���SN�+��Q��!*od�~���`��B��J� �NT퇅pG󌗟=�2U.~�W=��o&`#��;:����CeӁ
ʹ���{������I�t�+b��By+�(�xY��p������u���b�;���%ͩ�ţ�zr��p�.j�y������u��P���L���$�	[Td��"���Z�^Bo���^d�51n��k9S�~n�vW����wiD�PN\��8�i�;���Ӹ:����j+4��J�0�_z��W�{���S���J2�8N�##$�K{�^Rrآ��vT[�#�`�����Cp����Ċ~$�>� �	�W�o��˄7Q_� �9%@��"Ŀ�����IE��oe"�R�1�E����!s��ۨޭ�����1BS����G�ݽG���;��hi_T�-���w��5m�o���=wP�\q�
rm��-p��׊!,�=�&������  3�^*���R$�;l0Q �5[�F���&̐����2�4�Xd�8�uF��+�����zD�Ǡ�i�k���䘺(�L��H9�*���{Lv�d1�=�m<�'f�����^W0I���K��K^���|�����Aۤ.���Eg]�"-:A��6��_�A�M%_�gtx�vY0�|��(����l�o	pw񐐚� ��[T�u�z�Q7�V��5!fT�����x�r~�J�\Pn��l�Y/)Dk9�!����|Ü�u�|Ż����z"n�0B��*��4�^���v����ͳ�~0��3h.0����)K%�KF�luY��<�������Bz�{�2�h~Ēhd�h��ƽ�*]��V]��G����:��Y������
6�B5֭�i�J��F�D2��L�D<�W�v;+���-�
R�66���c�)�
9�;�=���1�l���O�7`\�D�.ՅF0%yw��;F�*������G��8�8�2Cʤ�I��(�,��bH�g�b�IP:D��L[�/����JX�����1����q�����'��\��N�O�iq�-c�r�/#�%��Խ"U���D5��x���6�tz~��S?��H�_1θ� �Q�YV]aa�4��e��{KG��A�^.;�/����+I��ʭd14t��lA�7�!
N���˄.�8xr�����VU�C��x v���|��[Ӊj�)��q�<���� �j���xMAp7E�L�F�7�l[�n)����k�!��b�8���T����rEg�po�(�;a�Yh�x-q;U�lQ�f@q��!�_�zu*����[CAjM��c �ޅBj�>��-w0!��'���=�Չ�Eg�WU��ą�dԅW"�p<���p�=ŀ�M
���.��>>��$����,!a�
��;ʟ��T0iG{���;��a�ٜ�)m��Y����PI=eA�(��NZs@~4v��_d8l�b���%\w�m��4�� 47x�{��xX?)�����+��+O�4�	���N��d�z?D�n�՛�9�}��`}wGBxs̫�\X/���j �)�)fKf�--gQ�@X~(��҄�$���x��^�᳉1�i�pc-W%�q�׻B!|�0ϻʔJ#]G�`�T��H鳌�?�B_����f����t��x��0Y�mI�1�C�T+��"�Oh��U�_���x��Ff+�������_-��+��1E[ŭ�`8�e#1	�L7L���Y��|��`"��|�]�1�������/�<h0�0�*���=ͅ�lU��ʲj:��>}q�J*)��Q�+���[�Ei�JbE{��3t��׍���ͺ��X��݈�����+��1���������JU*f-] |� �#a��Ɩ7�FB��m�lֺ��PY~i�U��.G.�.�X-3P݈�䒨h�����*c�?�}��z�� E�tءh|β2s���v�;�� q	?�\oq�7�J���+�<ϻ� ����{������s��e���p�+dCR���u�� �<,�R0pʦz>�\��|f�\-RϺW��y��_��Ws���8�/�i�9�ZnV�����T����ܮ�O�+�IZ���������+!ˉm�4vm	�?�FB�ז�%���ym�̙�h׶�t�ϐ��kַX����ڱJ^\���D�o�7�����E����Y�"I\m^�̦�e�-+#�D�i;Y�|�$��U�r2�Jɭ�x%\?�G��탒"�w�g�����Ċb~<w1�	�m`:��U�t�/@��ȲQ� da3Q����+[M$҉О��|���|IE�قImM���efo=v���YW�i
��T��X��\��P��Q
XI2�/U�k�Ѭ9�����~
��������f��aoAV7�g=틐p��c`�`ך��0ڙ�^�[�x�:O	4�R�g�5����P�j4����Q�x�K�������VcZ>�}�i��5x�Z���&y�Ej0h��/'E���ػM��<,�[��y�}�5�'��@��cu�W��={��Ksdŋ�x_�)cv��Vk���-���e;�臰zyĳ�dL�L���Jpy��ƶ6A-�h ٛj�khp�k?hC|��g��A0�3�v'E�n"��O�F:ě:�����Vсd��I.��\v�a�䵎���u�K_j>���w��3'WN�|O�@-�ߣ%�f�f���C���uh�R�"zI �ܞFAysΉc_��|���!_;�������7�2��	��Y�77���~+�wb}�IX�� N���##!�qAP���C�o�?.n�"��O�^�(r�#z����җu����b'�V�ٵ.D&���۰ֱ��K�r�0XW��`c/����,��B}#��%� �2�=Oh���)���F�h|��e���) un��������NbC�_+s5�o���b�tDb�PE���T�s΍X~c,W�fl���P2-1ޯP�	g�$�Rϝ�[�=搳���l�c�2�v���g!��*��D.	��Hs��B�#APK��')�fT�s���(�hG���\'R�˻����ԩl&��%����v��� g婞��{�s�����,�&��":׬�,!��֚��/�Jp15�{���(6�l���M�zcu8N#��~��:���y��?��]�`�v���u-Д��@���M֕<=us0w��S�M�vP=�|�Ũ,6�έl%7�����-O"�B6u���g~�\r���2���ڵ�����w���`D���	�tq���G��t*���&����]���Zi�F�ȕ�Vmw�"��@�,j c�é4��w9*����ą~!�����;��\�N�A7-�4]#��=���f����8�2ԓ�h�����O�9��)��m��n�%x+�l�\��-��H��}r_:L���}T�i���V�|A|5�����Z7�^�~��P�^��A��` -�3�~{-h���~KkU�3��}��a] 8���]ҷ�N�Oq��8�ҧ�0gމ4��`�~�B�9[����K.h���	fYw�pǱ_��(�/��i�X!�r~�YBq'���s.OP�e.ܼ���-�y"J��,U�y�,�ޗ$-)����?1�5A��*^��y�K�;5�����#���` �.R~-y��G-aCB�rm�]��[�.ys��Ͼ��D���#�����^[���3�d�c7B��+�J����|���TG��m:��I�?/	Ep�N�D�n�6?�_�ڤ
�~��hS%k7;o�ܷ@�x�!��n|[r��p��Z'�IQ�!�˚� ��3�uc������m
 ��t�~an̾����F��fA�ǘz6���������i�m��`�qU�яM�F�����Ep�^P����L7����_%ۢ(
����]�Vh[�4��:x�'�����3NW�D[������A#K�'�p��$����&տ̊���p���J��y�|��xŷW�:��^̽�JJ��b{�	�t[˧`cK5RDqI��!)���V@!�\)5`��6�������j���-W�}KVW�6`*��F�z�/��awI�����p�J~�ScnZ����c�B���#�C�Ю1(��
6��j�{��6h�=�#�O@^���^r����}WVȠ�.?�n�S���= "$��C��$�]deG��ן�L���l$.$Q�8��ʂ�6K���<{�[�d�ƣ6V�s�g/'�[��f�V�:	aay��p+�#�}:EL���x�t�-�i�=(���N�3�k���T8��R�f��y8DW�4�e,�3��pv��ͭ���U� u;I�W=<���j�j�w��A�����H4�PYEQ9��;a�C�#jb1�V�EsV?�)5�-����uRT�FOΑ�w-47}�o'M��~����hg����E����Ĳ&��eN�������;pZ �J�:�>����Eƞ���t#d9�&��[�ıU�)G�-�T��	���x�h|��D������Fx#]S��$ѿ~�L��ٝ��� )���h�}�w���� �'u��0���ǵ�+o��Nx�R���f�1���������rMX���L|������Ì���PV��-M�25u�dvu$M��њ� 9h̶BfܫtlM,�7������5����\�R�)���W��|�%bWeMe��?Yd����+	q��/���^Mo�ٙ���\�;Ufd����i����yڄ�gtf01�yq(W�m�KM�GC	٠�v����݋����[��3-��Q��Ϙ��h�7r,�3&��D��x_����=�����OC�eä%l�U�!v��+��؋�y�fW�cr�J�ƺ�t���}s��]?A�
7g��Zs�<�Hζ�jo�l�kZ|�3ט&�=z{���]]-��DRb��W��D>m�0��Jj���|$u�t$�����V�.�}���3�~�>#>�@?��Hg���Ľ�P�ܮ�3V�j���Qh���Ք�������x�K��]._�;��3�s�e�<*!�����}���Pl�������K/�m1�^=�A�?&N4�iN����1_/!8�e�L�m7x�k�0_�����k�kKB��M�S����.;ND���=�Q��O��hby&+E_����NI[�֏u�������/�i$7���~�BN��(zv�8ݜ�X5�9r[	h T���2_����h�Fu����^چ�L���~E �'���q��WI��Y3�
�ZL[X;c�"�e�Y�h-����A��G�*��}�ER{A@Z�o ��~��\L#��3,�x��j��a�ǼN����uNd�CQ���sT#)B.5����D�UsV�5b�n\�:�=n�����!�����P�hi��tub��Gcv�ܖ\Qô<�&�]��՞�Q�[����5�G\�	a�3�"�O2��i�W%T	рW�+��������O�/t���߇Bf=��B�9uA�RRT'�t�9��ڲ'~y�cl��I΂���0�g����07��>�;^5�%���e��in�3F�Eލ0U��� MY>��b��+4B�X�[P/�������"���v��d]r2�ѫ�ҩ4��E����7}�´K���_y	j�Z�^q��H�� ��`�pl��~ט撔�&0	�q��_A��U	��s�*!�����(�Ơr��ڻ������E6M�{O�^a:;�(���m�G���K'*�D� w����v��y�|�;���N�@�"��AK]�J��w��
���V?q��<y��J��uC�()��%)X�'�2[;.JI�3�i���Q��y��d�����!	R,c��:�S�w��+�з����"��8O~1Z}v�:͗�q功7~�b������)�v �B_�w���-���x&�w�5���hn/"�g�M����K�o��\:��Ɓ!��Rk� 
e����3��dਸ�.�w�.�P������C� 0�Da����ۂ[�3uO�K��C���<�"jȰ/�����Zұ(�5�%Rd]@t➷���P��J!�d��f������J�^ۂ�*?�U ���4��^��@��]��[L��뜓��[1��6\�͛�C='q� 7�m u��;A^n��9��JJ�?�Y���I���������S�W��K�?� �i��X���P�����Ѧ�ܶ��g'j���#�l���^7�u����y��@�Q�7��t�gSӋ��8\$�XaK�V���:���a� >l��Ȃ��W97���Dt׎w�Z	j�h�Wב�d0:ڣ#_Å�6�WUp������,��?�ܒ i�Wpk'��:9�������p�B� �����205${��j��<mו�W#�0�\l�RM�E�����;��/� ����j�ː}*���eԸX������A.�]�)��a�A�u�sb�7F�{��H����!`�K��� 8�#
i�R���Mn␋�������P��]�#�����_�+����N% ��6U��`
ɇL`�D.)9�p�8Aa�Q������:�a�"���Sp^�����vŋ��$��C�bԴ��q+��IʪP��:�M�ى�})��V�)t� �b������S�i��@ g�x�����\���F��w�j�����1?I�;ΆN
��]E��Zq!��w�M�EC/(/٭��p���J�aK�HVgx9����:�a��\d�d��_������(�u���L����9q)���r:�=���9��jn��m�U3���a��%���V]��U��-��̡)��q�
q�T�2?�0PJb��bJ�e��y[�,��R4�f�*���i.�O[F�S	 ��P�D�Yq�hJ��%��O
��Ԣ��	Kw�r�C��5��j�N���E�f���9C=A7SX,�?��� o]�0]؍��oʖ�$FG	vʪ1Һ�� (�.�m�w�ĒP?��Hhփy~
!�x
��h�EP�	8�U�� oc8�Jq�o~�SZ俌��=,�m�p��<�WS���lߕs���8��u���뱔�'�B;B�o�d�7D�Nr�VM�E�0������a�����
���r�Pu�R���M��� í=Ǌ��".�?=C�.a!c�T���4'zQ1�\�͌�S��w�ظ\ⶴ�a�ʐP�3 �&hY���[7�&�y�~�=i�֜Ef&����/ãxv ��5���)0gW��f�iJ�e�F�t����z����@�	Q8�V�w�y���E��������j�
� Z%:+;|�v���O���=\ɩcy�^��8��ss����z�i�0u���R�(��}��Á�p������i!�Tpd�xM�s�,Y���3 �(O!	��9N.��d�9GorX#��ċ���;M)r���i�f���r���2K�A�2�zCr�a�J�K����� �ᕿ��A��hrB���~�n�s���<I�J�3U�N�A+����%s�ͫ� >�Xk�6D��3į!�$8�5�A�-ߑ����1���	3b�g�$q�C����?�Z��d�V�T#��!�����k�r�Ea"��?����7�l�*�w�~����,O�u��B�i�M �X��#�PW����(s?�z?~�����&��f��9As��q!���*����G�qE��b��If��q��h
��26Qs���F�^&�>߬��p�	aj{3��v�ֹ��G����J�K��w�Z?�dO,���v�#\�P)⨟k9&��#ƿ������(U�!�V��;�n<�V�:��!8� R�}���?A�ɵ�P黼�$�!�1�Y�U�2ឧ���P��$u�V�a`>ڞ���h��v�����(�d^}��*�l�)4�L?��q+�7�g�c��hQs�2dv��Ǐ*+�!yo��ӏ5M^sϢ񡆣՟�(���)���B�t�9B�DO�pb���nn3j���&2��i�/q�.z�1�o�3��l%2���ǫ�9r*���.�}�ġ�ؚ�av�}Ѕ�
��\�>R\E� ¸�Ն�[q��>"<�K�{�8�f��tr�0+֦a�my�S�>^mG�̧#b���@ �W\?�B�������T:G��� x����N�h�`�������ȟ��Q���������=��C4,�B��R��:I`r4�m�kI�p�C��-����6�np>��]�\�ɶݖo2��a`��G���!4,�M���W ><>�C�i�UxY�%�g�7l
�٬�g�����F��啡.�u�8������T� �D��"�߯�����.�Ϧ@7���-�:�3DL�ҙ�ٸ���J���M��)�ձ��Ø�)1�BY�4�����)̟�^�y�	z(ǟ��I#����֚ɖV�-�� ��2�M~_'��<��	' �k�����P�V*��o���[b����R���ht��s�u_�P��?�zi�m�t2P��y=I�[�w?̵�$������}�����A�b�/^}"�Ky]�__���f�{m�!U�}�יFx�x�;d����� V}�Zh������i(� �+)�ąj��a���h�譭J��N|�
YV���S.�8֖�6OU��&^�98�'XS�Mt�x�3��v���75�ߐN.�3r��~�Ѝ3��+_�:dS��M�Y&�l��|�a_ˍ��z7���x�ON=\�ڴ<�k+mY]0�#<x����/�zv/H;��{�̿�mU��|����,|]�H�a�}G�J�2��<J�:c�@U�3�����e�0�$���7�����4d	�Z]i~�X���)ݣc�|��i��7&�N��Y����������Y�|(�	�C�~(K�I|��JCv?��Ŕ9G�}���z�fp i"��'�+�>����w��?����#*�{c4�R�v鎃ܿ����+��ZoP�&>�7�:85�@��>�:9w�䷪}�܍3h��"�J<�/��������E��l�ȼ}M����{M�I.�X�����kp��F<ҋ����r�����*�����G7� 4{P�f�z)U�k��W4�iP�ho���*[G�E;nj���rr�^g0��T�����=��a��ݟҤ��J��q)�b+φ��C!�R��G�GN�:�e���qH�#	�'�wD���DK����U����h�A:X^���hLҎdx�]�Y�P�^
.Y���1��R�_HY�?�{Y����/�WJA0�i�����6��2`�/2���{a��i]�b28+o�@�y���g�
��A�4lW��"n"��X7t7�+;�	�X��s	���M�9;q3,`h�A,��2�HHå1xp+��qr�Le|��E�Ѷ��{�/���<�S��mfDH�A�[�%�Ք��@��g����#�k���5�U�O<����X~� ��*�P~W�wd�t��y�����������7	��1޴��?��4��TY�~�����m�l�*�AWc뾚j.<�?�р�ە1h�p�����b��R�m/+�xS�R�Z�������uf(R�,����#uh�x�b�	s'��=GZ�t٦Y'�F1#`!�Ƣ�v}���>;!��?��?�J�������r�$�ߥ�"j�tk�����g��|Z��5�Lq�j�Ί��C�.݈1��ĝ��j�t��'l:��c���JӾE�҂�((�/u�"��6=� �w���N��4�A�1��G<s.KOK�� �4��J%c��P}$�Q��_��|v����&>
���V�
[Wb�3G�ӻZN-q(�`�ȉ�^M�M�ě�V5���!��6$>VG"��O������ݕ�«\,�mW9�AC~v(&�y��&S�-�A��b1K��@��Q�;%C�V��u�BzO1c��T��؜��Os�����׊P+ӗb��c�IG��4���ю��G��qeD���g�����#u�~��a߲��i9de���n2�C����خM�Α�ke=;g	�QT�#"�e����h(��~��U�h����E.�ŗf�TM�el���x@@�i!{��7���}Zq�Ȧ�]��"�|��fY����aL��#L��%��G��  T���#�	��I9�u/ѕ�ϋ�)CK"�G��4r�bG��tBh.v잃�>�~��{-!,U�a陂��ĉ4ՐDL8t��c�H2ب���8��:=|j����m���+�~-��"�!�?�+��DX#������`7��|d'�V�,���
>��4Y���Y��m<�K���X@�ψ�2�?ne����:w�ߐMs���3��,b�6Ϸ��D�;��v�bG�U{Q���
r�P�}m��eR�ˋ䶀z��O˶�/����b:��-R�L��Q,w#�*�uO��|���3��� ��%V:��$�~�CA���gw��$.��闞.��9��e�s%�Z��:*���(r���
�r�oQ���ֲ	���^݃�"~:I���������B�L}�<�c򹢂S1��w+&L��9m�g����!қ;r!ك%gA��(���j���S��'8��|2o�`������83�k��@ϧ|Z,��:#���j��nIr�u%Z0��1[�ɨ��XA{C�p�GhÏ	���_:1ß����G��X3�X~�z��&��)l[�M4��77�4У��� ��я�2��.^�U�PM{G*S�}73���!�$k��u����5|h �+��`������y*��u�6���z�PJG��DgW{M�F��Z!�x̨At#�r��mB��C�����jOBe���R~R�9eW;�"���ǅ�O�1��ĳ�L��z[��3@�0���q�OS���Y<�ڬ�Ub�ɚ����"�����u��;eu4l@"2&X^��8&�B$ �F�._��K�����kB�"���t�	T�+:e�pR.� ��l(���
��:�sT,�#n|m��t{���Uת�w5�lE"��ɥ���U��ᔖ����!���0��QeI��1ɜ{�L}��A�[Ʒb ��6L��YF����`����*{�סg�5���ob�Q�͹��,B����7���,nv��s�׋|�0�^NE��t(姶��'~��d��cRF���Ӓ�l��z��@����'��6�h'_��M��ݠڕ��X�Bʘb�b���z�ڧT��lI���yD&���� ���&��'y�Z�i7�I��wh��&�$����ba�:��������+d+9H ��GK�x�3�a�,Z��.� Q?������xl>k|�T�cz2RgU/����
���X�����@�[VN����&7mq��k]ܮ�9��5����m�l/�K9}��CI��J��8�_���?GW�y��QOH�UR4�^��W�"�#�Y��!�i7�ί�K�h>x�(--��y��Ӫ���n��z}	rV��1��l_������ɾ�8צ�F ��.X�&Gz_�Llu��0���܉^���-��*@�Vt�n��'J��c�������������p����K�����͠�Ps_.�7טЉPB󸊳�*�&��K���Xfs�~S���/�{���I]��k��ꔞ�Q�d#P���~G�I6�fY�ui�h�>\N�1�L4���☭�0�ʁ�����_̯5�Q m9o<^%��f|&����$�!ȪC�ʢ��&�-E�4�-א���8�|��7�L`c�br�R��l�&��"L�au����<��<��'U�Ԋ^5U]�%��)�)ǎw�f�{1X����L˧U��J��hKrJ7^Bҫ(�%�V��~"^9�wo�Ar�>d�hw�e�4S���:��
W-��٘5>?��x��%^�-$��;V�V��`F�h�����G�WN`(_s��1/u�C���$跈Y�;�����d��r�S�1g�!��'�U.](�4ϖA���a ���j�wy4D;��8=�O�͕�ׁA.3ÿ�%��:�2O���ƪ�ub�	��,�f�U����Z&d賆���n��ɱ�^�._�io���>?�n�숱~�airl,429?Vt����C������*��n=x��<s�$t�F<���w�#vk����@#0�F�@Ķ�*����\_�}�g���	�115��o�H�~K)���gjҧ��MXca�v/��f��ቚa��LHp����S�>@�C�����8��y�FM{xM�͢��W��ѐ{|l}�l$T�N�D��[��`[)�+;k�� �ī ���>�V�����tc��v�'�|H�(%�\�OUK�=�	����Ly?v��!|�=F���oSz�׭Y(��f�
F���F<�q�+ą��Ǥ���p|��԰^5]���^��m0�a�ގEl�s ���'�5�1����y���Ȳ�>Ё��8�f��<1�GP���d]%&UU�;��Vu@�U� ���<aO�U�����N]�z����i��n�ҫ�*�B5̓^ ���+�4�����Ѕ�����
oU���X	�a�6ElF�s��LB��Ԋt]T��.��0�E�o,l4��A3V�.H}�H3�/$kgŐ$:)������[�����Ĳã�
���}��G�D�A'��̎p熗3j�d��48h��@�gӛ]łI[c�j��f�r$J��cm`�#����:3yp|�R��T�˩�_��;���*��rɹ ϡt���p|Tb/�f}���H����3��z�K��6���}mgv���{ߎJ| \�uRk>��O�ıd�b%5�݀j�r���98g=����c4��d_�k_A|0)P��^Lr����ܦ���gW0�4���.��(y�E����h3�P�N*9.����]�gȓq�=���ؽ@d�u��
<�x�u��[�I�5������$mIO�;}A���a�s��X�>=��j���Xz�d�aS�Zh�a����7r,`�ʴp ��i��6��cr�Q��|+��\.:�����ΧKO^4����j���ܿ_H�1B"�OZzt�ʁ+C;��ba��͟�M�0)�E��H#h�3i���Բ�	�znV����-�&��:�����(]ɖ�κ�p�X}����W[�� �h�װ���^�֒�y����#�dr��A���&�����ʺS��l@O�\�IV�9X�l�	�O��x��B_�]FN�ށU��1�MQ��.��v�M��`�q#�����k��ݏ�Q3jB�����Ȕ���n���O�7��&��'���衟r&���$aR���R�����K�
��	��]��W�۶�E�!zCY?��z��p!8F&�R:BH:��II/��D�K�!�E]+�%�1���̷>�qC��˳�Hܑ뙽ޟ�X*i�d��U�6l�|����B4�&�J�qr���_�.�htX=_�� +�-[�g���}�e?�ʎ,��}Oid�� a�pC:�2�M+�-�/��q�*��n 6����-�oJ�eDI;p�Fuuم7a�,N��տ̀s{��sv��tf��aaU#����,�&������<X[�^B��M��C�W@��Ï�>c*6N�[u��E�$g���\�q�޽2PN���0%c���,:>�8�q�̅4�+�[�a>}��k����C��+x��8�GL�h���G�,����a]4�ٺ�qW5k\ ��[�������p�/�P��@��[�5�.<�D��6�G�k
��b��{a������טzE��ɚ���Ȉ�v�,R�n�1^�1�w�M3~�e��Ah��ʷ��n~U�����3F6�����}*�'��>C��~����62sn%т#"�C����4Eڕ��U�C�+���ʄߔ�sI@"��|�}�x���Չv{�E(�j���>"�	P;=�����"�w����1+��@]�xws�xnm�m�I�=��D?�[꾕�H�%i��V{�%ά���:%^"lCշ���ʰv������(�U��)�5�i�;�C�ڿ�Poe�TL'�����67,��7���2��k#���ED�O��O]��b>I��헧����z(e�(�|���(��Pgk+�\�"��xXs�e�xE���ϩ�x�oR
�2�Rw5�8��\�/�P��9�F��4;�2�`\�<���Qq�|���rX	�,+r�4���fG6cP�*������\�55O����k!���s��]�E����He��}Hq������(aI"����%0]<�!>D�"���N��8��ed�|�0�2�;�$�Smz��H~zȌBb��S�۱K5'�
R ����*�\���j� �B��7�٥n�[� լ�p��L�Dϋ���k�zr �Lا�:�B��t?jG>����,��3#p�b�X[g�ۉ�f�0�v�t���re�>3���Xy4�O�V����셒�/�����ݹZHe$�~y������ضP�ւ�d�a~ђ��\BT ��r�C�X�\x����qi���%���� Ḓ��k��@yF�����s����x+a�|�Y/Z+�� ����7�Uj?�fq�cJ�k�ѵ�S��U8��Pc����/z�}�c�AP��岸��\�O�+��^z�m�$o��6����#ʠ�*~ԇ�1����S0�
f]�n�(��~��ydp"�(��;r!�3Q��)�O��s3����h1�]R�3/��}�����>6�W)�4刬��hR8����Ag��b>[v�4�5�_{h�p�������!���	8������L)m=L���7ЇWҼ᭞������l��m��u(�9_ޣE�c� ��ql�S�f�D�K��U�V@�s�$�2�:�ŀOl����KI�k/�'���E�3��e�ۏ-{��~B�2��ɂ�jr��� �Z)��&P�A9����V׊v���,�n���#E0�'ǁ�<�E������`tÐ+mb��W�i��\���	
 ���_Pm*BAQ�yl��B�/?2�C`�c����GӋ���s��x�=+�ع��luP�Kʍ���:@0��D��&gV���+C�b5��u���sUO�U��<�ԡcnt%;ֿ;0g#3牞R�N��Iٶڗ�����'�z\�%`�:�"(0f#��x�c2��� �o��] �ia�3�?�8��p�O�u1i������I�ŧUґ�z<`T����Yi���5��oz�g�+�=���7�=�XG�Ǧq�����r���c.��S�a���6��Y1����Փ&v�1�R������CR���Ay�ѻra�mcX<_�^r;n�IDDL�;�DD�72�W��PE_���L2|���"J����&s������f(Bͩ�2�g�ѕ��������bG�z��A�{W�Ҷ���̪{�8��(�&����S`�xW�����COi�a�W�r����=ϑ��lZ
{��O���|uM~�Y_�lc߬'٦S���a'�M/A�3�Ȕ��N����<���,�l�v@Q�$j�U�el��Y���Yw_�՟l����7;?�H#���?�Z�[X��lôqPp�.���[B.��1|aH�n���X�7~�����M,5R�i ���ǘ�M}����О�@�̂�X�èȖqO7yc�]� 23�ٿ���N�+R9';�R���Y�>g%��!D��H�s��}3T�n>g�/ke�A�	1Ĭ�T�m唱�sUW�����IrPB�f�������h�x�S��G���L�*��u���a����he��-G�c��~;
n���F��:l( _�l��upfY�^�-����loS�����,ǻY�N,�	9!�.Y��(�{Ɋ8/I��nδ3�� ��T�ɴB�R�	ē��u�Q�X�>����U*9��DC��`h�Ԏ�f���l� jw/�U�ا�A���[.9�h��K|�9X'Z"B�������I!��Ƶ$���$��c�m
BɰˮAH��H�7��R�쁔P%!��Y��۹��E�A��)[���cM��	��V��6;R����bv�l�75�-8�)�>��.N2n37Y\cU����?�-t'�9�+	ϳ�XhkWy!K�~-�]�3�Fx���ni��z7���]�uŷ^ڗ���^-�"r�C�k��mX��ԊR-���<W���c��s���+�P;�\̓&v-z�eׄ��z#�=m��
7�Lx���!���:�Kʏ�
�bk�7Z�a�D��V�=�����X F���!]�c�f֜l(X���˦Q'��m|v�ơg}��cTt��/P������;\�a�?����d�p�/�s���q ��F���[f���β>��Ϸ�,�r��sL��R�<��Gk,T��4� Z��(�e�c���~��Xf*�\լ n?��-��1֮�͠rt6,S�:ڿ.��8(��k��<w&1o��3��,J�'��b��+�7
�
�^�wSB�����xK��t
�"X�ڧ䫩���fʚo4hf/��ڦ7+�5&d��4�D��f<�3�4�"�8��ۼ-���o�:g��= m���nd��d.Y�N[��(���	w�+���w�V������!+�7��;���L]-(Jfr;ʽ�ʽ��rD���p�g���h���w/5a �����ҥ׆\׳�I��U{�HbE�����#H����Z�_kd\��=��難��_�qK�c
hk!���Ϻ��{GQ@V�HX�Ҡ})3_m��h,�R����-G�@�r�V�Tsg�]�~�i�Gq�N���/R�KݖJqM����0%M,����4��� j/�fG���W���S�2��B���2@Mk���(����=!�6�/�fB_bW��ƌ#a�t����զ�ro���~��ݾ��F�_8��+r�!�`�Y&-9�\�1���9��(+PHt��߽b����Mc�}�D�c����⾉��
��/T�g9C��g�ԨO�Sɯ��|����̰��I0+[�̹$x�V��+��z� �v��v�OWnr ܢ��ء]b�X囁$��!�r�i��/瞋���4x�K���}���r����*�� �
��^T��R�����>�mfh��[�F�����M�V$�ᨽ���j�H�nKN��+`����4'-Ѣ��0
 �t/~��d5�JM9`�~�����M\((#Z���jdJ�$��#&�>�v���2vi|��{�n&�p������ ַ�V��5���'�k�pSdl2cn��T-�!�#��Օt�fy�X�4���e��8��X�n��V�Kw|{$���bOi�ՒX�"��iӷ�v1.>c��kM�\?ؐ�1{�����ֽ.��L���&n�,����*C���y�򬆐�j��������g�Q`�����B.8��������n[�E]yo�f�|���N�)D��h��ȉXWH(�~U��,9M��*/TU��%Z����y9�Q��گ�?uП�}��/�h���A��4��u�/��yNQ(0���.��F��#&[+1�6)
��^42GxEb5���P�3A��Fv����1#wVn�c���>7C�
�7�N��Hٝ(o���~yi��Giu��mr��b�I�x�ٍ��y�b����W�g2`�6���Q��1�w�cXm��>bS�C����nbl�E5s���|��KȁtGQ�X:�wl<X@�^�5�Acv�f�ɹݏ���S�]�6^�	��t#�;{a����_�[NK� ĩq�{���@���l�~��4g' V���NvĀF��X�E�D���G�Efc�2���u�����t/�<��s@^���
4�YM8͆P%�B��{I��O.�DX���M�����(Y���b4�	;[��O^�.}����C��%��"AMZ��[�6���S�lg���Z�,u����f4Y��K6v���"դFx����|kD�8�V8��n?7@{[ h�߆�d$��� �OC�����5��1���Z5���gzm�������U{�uﲼ]����@n1U>�)�r��{
5��o�j�ۄ�z����vTd�*�ݛ��{j��~f
5f#x�X{� ^���)cG��)K���Y_�)�'�'ט�i%֢��l��w
qH�3��2GĆ�^D���)��j0��-���iJ�$ԑ�]SID��%R��H &\jCEq��R*�'2�C볶{|�	*'k���˧YXK�����V_��ɖ�Q��XMS(�`�_]�0V_QzL�CFOIar�����+Ϋ���^߽�����{�gmh6�x�*�t��f�t��́�6��I�Ʉ1��SCE#y��?�˓r�у_ݍ���r�]LҲ�]Hq�$VT=9�@E��'����)���3eJ� �O)��N��A�|�ҏ��&B�7����x4ko�	�j:�k�[������X��I @wD�Y*]/��ȹ�h�T���/�w�bE���2:����_�q���f���$�^;^ii ������cJ�.��
cG��Gژ���B�C6�������6	!M%P�� ϥ'����ݝF1��v��X�g@���b�=�#�����c�0W�S^s(��@~8#{��86�����⥍�N�D܌ך��I�4�Lxh������}����1�~��i%ZQe)D��$yf'���F��DM���i7�+x��P�Ґ)=�Dx��T�PK����8�\x?U���捁�UE�p�B`tfP���{�����Y�]�{]�����pE3��N�R���ydV��cN�{!�;{��A9g��R8�.!�Kt��M=bO��T� �{%k���Þ���ņy���O�����hܺl4��Rg�S����Di�%�PrP������LW��mP3�l�m���qXF�=����E|;��ga��W�1 �ʇ����]tK"����!��!O�CKZl�[@g�F��v3)ꎙlx��-$2h8���M�,{�*7��1���%���g^��c�S�}�??z�d�� 2�>�C��=��Y\���M�=pWf����l���b\��p|�\R5=�}b�00�Em Y��!�1������(���������
�Wu���8��C/qR[��ӕ�Z`����9�Ӛn����l:���Txo�@��)d����q!�q�F�yw����{3}{^؏��~�ao���T�L�n���dZR�t�X��F�8�<�"}ڗ�>���
���W�̹���U���=Y�>�ِY�{���ك2|T� y;�gն�|�c{����F҇K4�*gOd\��w7�iif�l3���4�C�Í�h/pyj�b�t}�""�T1Py.�6�����층x� ��+� d0`�	�W�~�Ķzܧ�?v�h�ġ����� @�=X&�HtIY����m�*诣�[�b%�Dp,��0����FN>����3�lB�]<jpl�_vg�D̲t�S�<�»��>Uk��!�&`��j7LUqb;���J��1�#HBڳ!����rmW0�ײ_K�^�˺��	6/��A�56�h{ɜ�y�"rJ@^�"�����¹B�~�����k���i�./J�hl&5͹�˙<�$h�,�;=���u���2$�g(�p,e��[�_��$����������q��B)�����WUvn��<��&`�5���A�4)���8����_"r�I��ҕ�/aV��x��Io4��� �P"&͑;?��aV�B�l���K�_��J9,�Vl<ƥ�����ol�1.L�^O�rŅ��%uPhP�&9,�\���(�w��V
���[�UL��t��(��Å���"���3[m;Ƶ�M���K�NC�(J�m�"`�[��9<��XG�l����?��a7Ǐ�/���c�l+��u�� �l��k��k��#��R�fؽ%%���M����D�ޚ#߮�� #6�q�1�|�|�����i����rm_��m�%�P^<hcv�/
�qU�4W�Jj����n��s5���.O:@̦�ۢS����a��QPW(#����D}��]���|����T��T �\��m�<�$�:V-!�@H	-����2�u���
�r��|d��̼�k�GN_����B�V��n����.�f]���>�a��:�����nnreٽ7HH�O�)��X�8>��e�rc��(��xdX�M���<��>���Wp�׫+�_��L�g��ї�3~N��<�U��`��x��[�2rwhI@�%��&:��{�tOU��$B9J��tm�3}�
���t!Dk3}���1��nN��+!��t+o͑H����W���
.5�� }���fh�Dv������G�]x+4&�LC�4��Ҍ?�� 1S&+c 4#B�WR���B�`��N��^)Ϯ̸�2OLW~E��xO%wvI���D��h(lR8�ّ�V�c�F�����H��`F�p����`��{��n��0�P�TJ�}'=p��*�d{N�6�p#C�h{-��b�P
[	3�}�wnh��JT"ф�_=pH*Ʈz;�����H�k=hӱCˎ\���
i�g����<6="%
���4��9ο���O3c��^�B���;,���9��f�������=�u�Ӆ���$;�W�A@7�?/ �֔�D��ia���E�%��/���<�1���p}Ƙ�H��5*���N�O;	@��dB|,qC�1����(�������}I�+ɵ�Ɩ�u|�$Y׵'�~�b0������E��=�@t�g�迍�zV�\9�%��0�wT}J)H�3�;SJ/�i��-��b�y�7c��B�"��S_T&��!�����K��}|�t����U������Y���z�-�/X!I�:Q�?����]ԋ�Z�y90��+8O�̵Ϣc#ς�3�|��NP'1�3����A��q^r�^n�gX�J��cR8���	&'|"�j.j�6]B�m���E���uD��e	��:�Z�&�1ޒ�?D=r�=���������I��� ���+�����aAڈ��c�
�܊�'�\*t�� ���j,�S,�4�:�F>ꡚ�����܁"H��&��4S��X7us�I�wg�em{y@����~�G�0,zsDڊ������Be�0�	4�XLw�1�����e�N�W��= 2��t��P���<�l;��Pd��a��2�|�+|��C�y�|(�ε���h@��A*� k�m�:J����ɲ�Wa����N�ku	��҉����p��a`k��)�kza��$�ʡ�|�@\��� x��^>){ck7�߈]{��&"�H���,h(B&���
dG$=xԚ���(a�#3o.-�����n!&ڣ��s���W���c-*1|m$+*w�,O�n�Z'&��ku���K�y�j7m���v��~D�^�ˀ%;I%Ge�v�2�P<�0+�@��	�����7��ȿM0����a�S�#�L��J#�����e��6�L��Sd�����q�_�;�_$M�)K ?ӏ��2G���P��E���-��<����R�H���B,�E�<-A3�������$����f��"��1���Y6��b�9h�UWq�����!H]
�׽�
���`�ɬ�u���ߩ�D4�u^��z>�5��:t�(��jud������
��iN5�kl�vI�m+4�5��ǇdQ2; -*@K(>�z�����ӊ����h$�B��~w�uH�� ���Ƒ�Qӓ �ܑ��ڮ�Lʝ�Wz���z��+*ԇ�B���Nе�)���K4c`��q^����-pM�a#�%,Ty%��uψWv�i-Q�K�d�3**\��IY`t����M����l/�m R*Y�����{� \�H��:&������.�F;=`�w��Y��=S���;''����|!+�@�!U)�I�Yz|>�=��u?D��DH�q�8�Յ�D������|D��bU�l��6-��1�#L�3-�Ӄ�=�h�1�����V�-�����/�ﶍ��Ӕ6�C��~97#I/�'m�X�}Ԯna�Z1S$:~����e��1#�mU�(Iv��W:����/*��=M�3��D�گ��E_'�_�¹�WWԾ�M~;��udT"�"OT(5ɇI9�Q��S����ʬs��V����i���Ŋ,�Rܗ�a���P�F������2�/��#s�¤��*������za���z��Bڜ�x���9ܨ��ܑ�*��"���/N���W�U䅇](�xlwi�]�?��D��x['��WQI���=�7�M�Mՠ�}�Fm�t��&���O-]X���7-�v����(2�}�H�g�f1&�}ʁ�MK���lU�Gj� ���&n�/�s�I�n�l׻�mAc?@y�g1�h���̉ƨkÉӻ�H80�M). x�*+����@��M�����?�~�|Y�x~1_�@yp���Y�ICY�U�	>>�p�x˵w==���)3t�Dȋ�ý"��W����;!Q�楏 .Ԣ�al�CP�˚����(!>�����D6�5��@����	�!���n����'7�-�<M��9ts�_X�_�49Ua���F�Vs��&�T@����LkA
�&�e�H6VA�cD�Gb��ʷ�@�rb��
vy��!:������]q�J��a�	�Pv
<q� �A���F�n��"���:J\�1�փ1S�Ha����(Z_��7��5u���� \�{Jfp��Q�N�����Q������<���ۊ.�>%�q¼�Fg���.g�T�Z�'��0~�����-9�*�fo�m�E}IOw��Ew���Z���Gi'9������6i{3�qr|�v�������1�M�3�0���ɻ����콅ˈ֖6S��WA�C�5Kv!����;|�E,y�a��1-$J1?�.��]���S*�}�Ԃ�hyF9��G%"��	
�|��m6�:�O%K��P���i��ƨup�D�̧*�����ЁXl8��m��1Lt+�V����u�U`�M�W�	ժ�O�v9�mh>$������o(�߬'LL}L!ߺE�� ZU!��s��\�q�Qد�L���sjrq�cn���i�T��5(q=�-���N�!�@��q�v����Qb�ɂ&��
��UeKU3�Y�ޢlՕ��$�QE0����I�SRH�v^#���xN^�0���2���`Ã�s����Y9����l�����K��$��|��9��?56u�:B��흔�Q�Q� >���w釋��?�<�R��i.uh�f�e�7��q�$��G��u*�����Q�#�a/7N�}�{�%W�)�[Y*� |	h�ǭ!�B�칳iJ'�]�d�0�Gs�\���t��b/�/���2�U�W���!�$�yr=f�[8���vZ��ypk���OP�5S������j�A�9���������Ưz�����ޚN�<t��<�,���-^�O�����2���׽�'�=�K�׳��NxJ�j��L���&���*��}�Rē��B̪������@9��m��z�b:U搧W��D=��%e����w���p;���{uQ�c*g�6��P0p�Er�4)�v}�@mn|�̇Ya����������{:z��-D`�J
�#�JvUs0^4Th6�1���B����=`H6h���Ө�Z�� _͚��-`��,�HF�|��b����E�� ���:�X+t,����H�V\��T|ԡ�&v��<D�7��A��X�|��%����7�RK²53����؞�0B�!���M����J��ҟ;a*��x�ɞ�׋,;"9z2��=�3��?�y������yƅ;9�Y�ed=&��_T�B<�t��5�Ed�����X��6ε������mC�3��M�9���ҝ���tDm\}����J�'�:@'H��Uc�x�)�����U��U�)X;��b��|ˌ��1u�R�qa��#��8i�[��8��N#��ܮ�V�H8���K��sh�v���R��4�~F{�Q6?�����a���	�'NE���G��K��/��\ȶ')�͘ݖP �Զ8s�`H�������$V�R8i�ۘw�y�w�k`�"�{<k�	q$�^9��x�-%}H/�1x��<�/Ӆq��d�8D^m���~��`��P��w���r�z�e�y�&��x��и�J�d
pp��P�a���^]	F�{�i6G{�%w3HVfT�F�mE=!U��0֖@����CgͭTm��B��3��n�+��l
���LÑ���Y�/cm��ٷ�Ӱ"�۝ߴ���{D��0g�o��R�o����F_d�f ��7�%��Ŷ�}�p�PB�I��bDo��U C]T�SL�s�A^��D=�o(.�@TI�Ӎq�~�:w!���?+�;�k�>"EgK��Y��Y�oC->�X�����;X��DR�%��h����6�~�׾`%*��ii�e��X�_�e�xx�9�2��տś���jU��'Ь�)xN�����U\��!q��H�yۗ���KhNд�j��FW�q������=��`�Ұd��9��%~����Z�zD��I�~ϥ�՚����>*��_#]�:�X]i	�-���(C�>EZ�8b�x��qQ���n�Z�R՛�>Pg,���s���ol+�W��?tY��Vfʧ޾-�ޜb�nO��S�[�E�D��HI�籘�A	9ޑ���3ˇX���ъjO~`K�=�?R�ly���g���'���3[�� �ҭU�o�(Z��kN��q��4�D��<,2qA���2���b��91<��Cbq ����iP�CM��yt1-��qc,�%��&
��)ؔ���`�Β�x������z5'R��'��wh���ZY�,P?�2Q�!��&�=��#��?��$���Rw7�����Tn��ё���D��2Ռ#��Tэ-,t�7"���KA�w==]�[�θ�H��_@����	�d.�z:G���M����i&$YLvl��`��rpY�[&���6���I͙X�L�0f�`2���ӛ
�u�t)!I1$�}���ɝ辽J�\�j�;@f{/� W��%ܨzʺ
�[N�vEM0�<�~�g�e����۠���Z���������#�t����(\��Ͻڏ����� 2|��
���^��U�z(�N�:��6p��04�#W���]Qm�7�	5���S�.����dh�~x�)��<"�o+�m�
pfAt~)q�tĤ�kA���C_;�%F�1�2f\8H�z��7;pEi��f�S�g�3k��=}�l�~����>eA��M����
����D.&��K!=r��'���>�}�c�k>����݁�-thVQ��@��e�ɲ%��9X���e���h/�[� Im=Z/����^�����7��y|���鮡���p�R�#l;��p
��l\�Q��c�k��(z����*�O(/s������,N���T>&;Br�H���Y�`.�W�WwW	k����l'�����o%�}��B�NGa������z��a��J����� �~"Ȗ��ɹ�i{In��9FQ8H����P�Co�h����8{���`�yzA�sf�+<���$�'��2�m}��N^���Qz�g�V'�����hT1��O�ɌҸ�.Y�A2N�n�>�M����ZS�+uI4�hRh��� ���Je1`S�BJ�v{6�5�r�h��aa"�u�Jd���) �;w�q[̝K��z[���h�(�i�@��{Ch��-��_�=�L�>�?FQ�]O�s���p�˺fdvk%���LV������Rꐜ~�]�z#*�<�G�,Ż����9]}�L�8^�"	��}����Pm�o�V@���ϊL`-��t3�W�����$Iq��*�dt���[l���zR#�ث�ɐ^��J�Q����~"q��x]��%�a�d����][t�����9Z_�A�7�#蚇~X7���4�kl�j�"��Wʫƈg�#rQ���;�k��Ϸm�V�rX�������xZ
��;�]j=�ڢ�5ҏ�AD�tgAv_]����уq7�\�d`P���2Ƚ���"q =�.`0}�?�E��Ï�G�P	ۆ����x�>��D���RX]o#i�ʐGV/NC	nf�&�`n5�Ay��������-��Fr��-�%���)�s�MV��a�OQ|���� �����D��0GV�p#_���0UO���ӱ4U (p�bb��ǧ�ΟK1���NdXK��@���O#�i�Ps�u��{�����J��_'�)8��a�:��(���o��ђ�ƾf��к.x:Q �^��f�[^%$r��0j��yor.�t\L����ЂHV�q���*r�b3�|�9�p)bZ;p��F��3��!�s�Q�Z&�[f���z�x�X���_��,�~;6��ϯ�zp�[��ׅ��۶��0Qn߬�\�`.��y�\�	��c�\ ������P�4S���"��� �lըNw`@?F8�t�@�:!ǳ�|��γ4��H� ���;y0�9�1Gz�m�,P����F ��j��P8=�j���9���0�(|XɆ����y\m��"|�"nrTڪ[3S��J�(P�I��xr-�^S�ޟ�2<@!]qı�c _$�|a	5�� �Q�"�}�m��^����ay Y=�x�jEp�c	���%m-8�kn-k���� �T?2$o�8#�&6c�� �,N8��ᔮ%�`#1�� V�Y�E�A��zZ'�r��4&���z,�A��	�������D�1� 5r�#C����F��eNAn�H�������|Vma_'�JѠ��ȋ?���/���i\��Q�_����9�)`t61�A~)�X���`�$��iɁ/�O�x��_�NӋ&��,?�u&*=Q-�Z5=�^���i4���(2�(D.n-���Q�wPO~�oԝa_��䋩����:d �tl3�u��c��[�O�.a����V�4I�B+��M3-Z+
$RY��D+NU�5��ݓ���O�dOfQ!3bon���C���*Y�����Wl:���V1�����p��+
�a&�t/�Z�y���r,����c%b�X�U���D���W��=a4uxc �}�bM�hq��J�J�����W�bzKl��+����zb*�~i�0r:�A�OV3?ꂤ˯�E�3����x�B
hA���/��H�u�!aoux�+��O��qs�+h���0���4� ��;�ps����F�*ź�#��T*g5�C����*���������j)�>�!����"��!I�禘e֢�(�� ���m>��Y�k~@��q��B|N���f-��i�͵\�����;����N�L�i�=zte���AA�(��o�S����9Ł�er�X͏CU;��jXj스�3���{E��I*����Kd�V���IE;�"w�49�*\w�SԻJ����gs3�/<^�)����Xg�:j�"���<sH����U@M��o�%f��8Z\�nj,��R51旅:�F�˗z�J{n���Q�95�&ш�.f��h+})��#����M$44�&+���R�$t�2�VS�@(|�g�D���>�ޅ�/ә����P��gOw�T)������š�;����ڽ���o~�n�X�I��Σ���
`�>'��#%_I��uXUĸ-�j�Tf�_�!�r?�͚�}��M�� �������B�T?l�����ǅ1�\4W�m��"d�	�Ћ�\�&��=��-�xo}��[E�ĘW
ءZڒ�Q���HTЋ:.V���0�ZU�7T�ǐ��!�C��2s����ջ��[�G�<�e*k�+%�����q�C�#�]$qq˛+�Q���d����e�v4�\��=�j�0�5zUy�j$�Ur��h�[�[]'�ZO�2Ѳ���������X��%W���[�"��d��Gs�-b�eď�]�}s�A���gr�M��\{sQ�y+��5^ـs5��=�RI\��&^�i��m����#^�%�h�	�Ҳ���!@����.E����-J 0q27s%T�4;�Ϋ����ID�~���x��}�`9���DM}�Y�T �Lc��'�#��p�q����g�Vt�C
�MAJ�0'�/04Z���d�*��G&��ä���%�>���a+�`���LD}{e�>p=.�'�K�����vrY�����~ΏR�0$�
-l�<:a�YI@L���"n�*�B�zZ��^�ek�5GU	hc>�F R���|�G�W��P~Ò�1��hci��v)f�Cr�y_"�O�q�ae :�@R�<G2,ʹLD��w?.�r0�ca��r���n��Β�㚱��_�7ʮ
W`p)��ZP,B�n]z�Q�򡡨'�˹HJJ�!�fr-�K�ŻĲ�Ω݉���[�49j�hc�sPB�e�|шZ��C+���%ui>�`�=�#�"joAS��;]�p��L�������q ^�|ȻM2��~��<��욄Q�{�9�I0�I���=I6��8Q�8!PrI���R&�r��htwB �8��k��_�����7�O������?P���pz�v5�F�h���.���͵��������Y����%T��O�.�v���v��lH�h��[d�W���m�N��̆��sH�|�V1 �m�"���P��Jl%7�Nk6�R�+��6�A��7>���{����,~D�e���>� 6m2�x�M.�u�p�,�E/�i5�+'K�6�X�ܮQc�g�#]X򸾁h�a�(yI�6�	�VMh�q��4������4���v����4�I�4vm��(��O_�Р<R�vn*F�^�lJ�n�uྖ�쎺!�n�7K�0&qgz�z��s������s*�y�������Y��Art`1�z �S��	B0��c�B��X�����$�M�k���yv�nг�ʓ���r5��>i�3�\u+v���ˌ�7ia_j�E;���c%��C�h0z>����լ)��śQ������R�� A{I�7�~H]Dn�֋�M׀n��3nN�a,o���Xԑ�#�m4�f)`�S�"rF+�kgU�KPu�Ө����Ux���$ֻ�n�L`$�#V�K;c�i �}�T^��������$-|�,�1��XJ��ײG��������+�@����J_�B�4/~s�RR2eJp3`Q��UO��C�D*����["3�Yg�?�o�V;�5�����M�{,������F`��Ԫ$�����}zXߩʉs��];�.@�S٤�����N�o��}0���:2L/�~J�۲���Qi�R���W��WG%<�oo����KBF"x�v�-
�o��6�L�}S���ws+��酘��XUp�3�Ƕc`�����X�5A���`�w����Ù��B�m.7��
�ρ;�*�$^�<"N���X6~>N��S�z}�N��R��c����/)T+x����}�$���s�Y��"��3�P���SD	�j��M���kGG0�uP��{\�R8hd�����v�7���!�ap\U$NV�õ��Ie�Q
�Y��k��W]X� '����E��x&(�����S���+�M�'�����P�����5r��y���@��%'j�Nv&?ͺ��/G/��E���=e�߰���V�DH2Wۈ�y�3WCx���g"`?@Swܿ|A�$���6���=sG��Y2�6�{Q�a�ө?�/��6�ܵ�X��X?��x�_��YSz.��6xJ�_Oԣ��"�h�F-�L$q׮9�)9J��������BK��v�(Ө����-/��ӎ#��?CY��>�O����2��)�|�X��c̀�,.�D��mq�!V1�㰄���@�o�T��vZ�*�U2a7�OL_^6f���uo�����i��2Cn���!�>#�j;�U����1���x
��W��1��M|�h�����l���Amկ4?y����V�����U�S:���mf)��`9��hT�>�g���xq���]r�	,4?נϠ ��
iZ�1�4&�C���۹��\�'��n�ª4�:{)�o�Ⱥ!��U��_Pw��/���Dm�d��`��>�|�����T�D��HZ8dC��\���Z�}�?c�e�:W%n�B��%�E����yJ���=QoZ�	�� 8��V&O��$������+�\iG��<��m]�  ԃ+�^�̩΍\_P��ӛ¦L9ǟF����L7ZRAm:��W�=�h;q�⸘�Fln�/�������)���ߗ
��b<�)�2�,R�<V�հQA�3>��6b[��#� q���z>6)�����O�rq��7��^Nz�B���eD���ru��㔀��2%�̸�[u�Q��pÜ���7}~L��b]5�U=�#��	�E�ͦ�f��k��Nf>w-� �$a���bU��I�ϭu_~)��˝��/8"��?h���Ad�V��+�x��<~lS�;p�q�L`���3��W<��
���g�2ѶȺ<�S���;fnI�c�xU� ���U!�i�� �fŴ�w��@��f�: ^Q�/�Ƞ{utIqf�����W�Է�F�"��3,Q�jg냤'C̙2��WP�����&�su�N��$4Zƭ\5p�x��F�*���q�8{+�t����<E��~���%U��f*��b�6Q�N��PI>mᇏ6���T{�Y-Z�s�N�N�d�)Y�yF?͢
���]�c��`<h(��} �` �4�}?d�M����������N,}u�J]�k�I<.k�7j��Gc7�?`bk��58;���꟞�Iέ�����>у�lK��QO���~w��b7MraN�St�X9��|b����@U�j4�0D�ڪ���RN^��<4�����m���Q$���:���^;�������٨�m�����A�\%��rI�F%T �%�|�/]��"��OY�b�͡ɿM��	�t��L�$ou Or�Z��R�jF�>`V�-�X5�;\�-"{�&c�z%�<�xg)�Y��E�{
�~=K������<)?h�SVO�_�ilx�CoV?��p{�sf� )���A\�߁�Ʒ�a��GHrj	�i�:����,�H:���:���㻆Ui��@��)�Yc a������h�)����!p�`d>�G�s�Q��If�gf2��5<l��=G��h��s�'s!Qz��y�	�ތ��:;�~����|�c"�1�|`��hR�?�7؇i~�/)��i��Pk�Z���dڱ�����ʂ��q �a�7���*�j�lByP�͹����S$CZY���~/���<�#e e9H�\��w�����+M ����k�/�<��s-���ĺ����[V��-B�O�zf�������-��H�c�h�Hǟ�sh�_/�T�D��E$��O#���,gL	*�[�)��(Sc�F�rHĥ��&��Kz�'�P�wc��а?�Œ�j�|����]v5tbc,y�]��D���@T��J�}��(��v1�ٯ|G���+J�I�F/<L)�V��+��R��9R�u���TԝbT��_OM0۝S��jEBr~Ѯ�������k���4��Paõ�ݟo0�zyK��O��6�ë|�LI���q�Y���<'L��_D5��)'`f��Bd��3xlꇭF�Ei�7�T]�\%��C�	C�<ܩTCP�P-��ͳK�y�r%�Xm�q\�Q�K�M;�q# �b�o[�Ȩ�����*��E����V�z�Hz�:�2WQ��:�wL��}��C-1�@/��uu[]����&�A�G�`�|ˮ�_?g&��x"Il�3��z�+��I���u[4MU�*�+�����h��Fy���l|>��Ӟt������������^��K=o�b�h,�o�x�s<Qi�1}dq]<���LS�z��"*��v�O_G���}S��~i��j����,�\�6�C63� �����dzD} ꆀ~:�R  �#U��$3��ʆ�F�R�B��+�fZ��C*=����ٰ�鴲?J$B*%����ʥ��3\ٓ�6k�Z�Y߼;V��=^Fx���-�0���|J'�aڭ`j���o�a�e;�����Ȭ4�$��v*��-uRE
�#{5[n��>�l�(�$6V7V*�<��$2��I `�\w[��Fi.�S
�I_E0�����b+����e������à����H܃|�D1;�>��6�(�ՙQ�?���<�t`L)e�^�zA
'O;��	�=�wF�,��D�&
xm9�۾�:ZX�Bi����,�-qAk*/� �v�:|���鴣��Yt�>�6���H�@>�4�O�Q~TܾE��CW�*G�$J�m�0�|�#(�Ex>2��xk���:�ɜ�O�]F�!��FXJ7U�F�E����e�)���S'Q<#G���{���O�Y��-%7=e���Rn��<p�x(]u�13 ��)����W�$Es��1���F�G��!#�3h���a+%��=Řߪ�oyUцo�����ɛ�V%�fx��P$?���n��h��ª;p(�C+�����/3�ξ�څ�c��N�%ԣ`?��p`'�o�]�.!�޺��3�߯�ƞk�=�>��%\g��C���$M��3�;i�c%2K��s+���2yC��S�ѯW6��7����~!_��fC�w�1�X���?�� ��H>1O�h�˰�Br�QP-�zZ��A�i��my��l�0K,����b���ҵ���+
\F�A\-F'�z�m�:D��qcEz�*|��+ź56���?I�] |�$�w�i��JF|c_�$-�u)�|�Ls���=<�r&v; Nn�t�~U`���^m]��  �=>��Gh�A�0����{�0|c�K���Z��p
K�zcwU��)}Y�7��ge-	-�wGS�������ܫ|CI��!��[�9|�Np�$M�3�)���mG�~A=�,F��Seo�,ba�˰�C�{QE!������K,&���CY6�>f�B���@!*��G��v�ZK��J0�Ig��EO?����Ԋ���*<�6�@TG�����;�c7��fэ	��A>�J���$�݌?'Q�e�Y��ov`9�"�|��c|,٬���#�䱋ط�f��}��ep��~O�tV=%��t;J�.���Y��5/������c�V]�Z�۷k'!�u�\vW�b�LwʴC����V��y�����VJeA�c>j�ckJ#�b��۾���~�aWɡ��y�~��3Y'�d{X�����_��f�@��5o�X�,���?�ASb}������6E���͟6(�G8DZ�L]��_���5X�^��f���|�1���φ�R%�urH��C4�����G��!��c6�����Vw8M�Ѳ~�JUh}�)�w�dT�x���a=ˈ�A���z7[����In2�aSm2ۓХH����E����Rm��r`��c�#-��7�4뼑�TH�Q:
�w��K�b��t���ĕ�K�C�=uс&e�A�y��h���s͂_���ҥ�[|]��zh{�|��#�F\7���o�Fe|oT�R9OQm,�%ϰ7�3�\� c��6~�]�Y���Ķ�����U�=����$�;g�Q��A0J��͗�?c�hxQX�U&�����V�Z�wN�ϟ�W,�L����\�JD�E�J�!�P��	
�Y� �$�ұ_�@ǖ�q�!�$�t�\5�nD�N��^�A��L;L�8z]�#iY~��^\!��);�E�8\�`���j������^���,w���s�LC~��*��FJ8&�[Gj>�����*.h��~��e}���,`���fi�w����{Ra���3��4�ӨI��)��	Wb�6\_��p?H����> :����P���ǶT2�ӡ�-Ŏ�8wq��n�r|�VUCX�;���0.� ]��L�T�CyX��77_(�o��b-1��N����e-��̂��>������^�.����C����@p<ѯ���!�1�N��S�Vc�x�n�V��x#�҅�_ R��V2�����4��/��w�h��|�+��-�����{��I����1{��������/|���q�;Jx����V�ס�Lg��`4��{6������n2���q-JaoYA����qH��Is���p�Ҽ��=�������C����$Z�Q��*@�kkR�k����Z�	t�z=[���qȝ�Ljw��G��4����y%L2=
�.Z�wD�ڈ~A�m����(^��R��Q,����L��ma���]��;@Q���,��$���e�6�o4�a������؝���3�b�W��Oy����s[�84g�<!�UBR>|��9MM.��W��IŲCJ2i?�hI��ud�c4�x��X���{Ej�Y��ٺv�����-�^߻���P	�soPco�G��<�=U=Y�����ٙ�P�*P�k��6O��NO*\Օ�01��douv�Ѯ��!O�>�D��CeN���
S�!��g���骞\c�+~SE��s��.�yB���hT�	�:L��0).-��V�e��o���3�i�PӕY���9��]���X��۔m��$������DXt�Q,=9Wh�&���S��f����e(ز٧�)��9�_P��_�@hA�F�˰F"�i�8��)�G,��W����QB�D#��ķׅ�2�	��X��B���W�&b��~ʎa��G�/C�-��$��o��Q+��du��iw�JÊ�}eȦ��`;�C?}Ƭ�2��c��{���L�W��-��{���;y��0�V�S	ٽ����Q�	n��\�YQeeQk�6�lo?�#�kb�̪k�L1��A�-�0��B�&*n���n��N~K��������|����ZZmt���(�{;hK.p��q���5%��O^)�1F����	�-���B��{�=�R6_���
�H��&�oM�|��{�Jp3�
r5��HltU�,!�kI$��a��"7����Aio��ޥ~h1'-ƈ��Z�>���*ԐL�S�B`�c#���)��wJ�J�2AT"����������s%�����_���W�Q����Ѳ(_����o%O�_����>�L,"U�9� Җ�������p��"$�j��9Z7��^6����+}d�W~%a)$I~����-mIdwʔ��fd�j��V�-���� �v>`e��d������|p��,Ǩ�� ܐ�����^Yx�R�{� U�:l�5h5�p� C��x��w���Y8��{!�sk7�D��QH�����Ǉ=U����|�h�H)�n�+k.��=�r_}�W.ރ�P=��}PMX��'lHz<-��P���j��O����3���x]�D�Ӛ������K-��D��(F�[ui	5�du��_Ē���(a���K��X.]oBY�����Q?�N��ۊ�Ӎj�f���*��_y�{$Ki���ߵ��k�LI�p�Ո�/�Z���&��[����d����3�+q�BQ�Rk�;�UՆ��LB�hì���� �z��$�SR˜�Hk�M� �m �����po�����0���9@[3_P����@�yOM�e���t��K���Z 0H�y�JY/�y�wo�h:�$S��<O�n�wD��`�� z,Ab��8^Ɂ�5a@�����q�����{�ʸ��(PTyF>�3N-��{�wq�c�}w9rqk��\��4;7��~����l��������E'Ry� ��G�r	�;����ٌ��6�9��V�s�����45��~;6��$���l�"�-^�)7)p	���
�u��oT)�˼�b�([w�f�>�@���4��eCj���w�rCp� �H��6���٘y�E ����"%��q"����c�� k�}��xz$��x4�}����0 �l��-�d�*-���LWen�qP�W0�/��c�o/�$t��݊�����^2�9�8�h���D�?t��k˕e��P?ņ2��p1��X�i�6ƭ�[�n��ԓ�ؿ���Ѕ�i���
:�1��Q���|��5�%X�����!g���#PZ�{I�ҨN����g$_�`E&�ߚuIz��hf�������E���XH��%6�zO�u�� ��T|jͰ���q��HO�fr�n�u���_��ܽ_�Y��2H^d^�������_xh�.������ީ$/��޷�|I�ub�Sqg_
��9 N���inf�A&?>a���MƬ��ժ=�T>�B�8�9��(�N��16f�UHO�`�9|C� b���h��B�[���;�-1_�]$w���~\���k�=-1�w'���ڿ ���w��R�����Bya���a�a�y��4-<�8!�N���8P��3��߿��3iz�11	!�ԤP9���$ꝇ�a��捭�ȱ�l���v�Z=���X��[�⬂�7jO�n�KӒ�o�T6]��E(]D�и�{pˌ�`�!���\6�)�.�ɖ�A_��b4�d������R_�S�����L{J�ǭP�H��z�������fu�+
JX����4�O�q���Z��[�-X(���]��^�g7���J�R��m����_W���s�Y�		�:�ȣ@<�%����Z��+�N00l���L��P��)Fk���Z%�r�Io��!�7�%��|b�}<����n3���Q����o����j��	�^�x�[!��E�Q9���t�qk9���&�Y�r�߅1�WB�W������I�ظ-�:�[q�0g���P�Op����=�pn��%��!��Cp��i����Ē�\ Q'5V�iq��o���K�>�e��pJ`M��L��4�n<�:'���˞qZ )�ib��)?r8��/�*�Zi�!���Eg��
R�,
��C�O9{����+3ZU^Z�Hi�����kہ!*��k]��2F����}��m�i'��@�zq��s��}�'�]׼�$��M��y�i�j$�\���e	��e��ˇ7;N���E��1�	��}�=���M���`O�&2��Ǩ�I��i��^�D@Z`�M@�G�����7�F�ۀ��zq��U�DQ���h-����P�B�hJ���:��p֮�kNm�G���.R�ְs G{ʔtF�n2��<G�!`����O�{ΔB�Eiwe�8�>XN�?��YԚ��ҽ%�ʯ�-!�#������v��a�.�}2e*"�Z��!9셴-�cY�ݰ�/O:u��*�DzRi%�2�d��H�.��
��^4�6�Ec?�K��Ul�����ł�`����Ċ^��l�.iG}[3u�>~��@�{/YP��������f����%|+�儴W$���� g����}��X{È(6���e	vn$�_�5��\�x)}ߔ�B�2��%/�7�9�������q#����U�y����ѠW���7n�H@�x���T3�@ry��ڈ��@�F�
b�PՉ�����D��
���zaO2/e��>�8�J}��vMJ�Jp(=�Ґz�� �y/0	'<F�M���$h���c��$�,�v�"���pv���'����eǦ�Y�i�h_�~g9s�'�W�[�6D�ט��&�T��(�u�F�#�	�@zbZ�gي������uBp+������-p��od&�1�焆;]a�a�ܘ-���e�$��t��zŮMܝ4#Q�K铚魭������ w� $��c�h������ '�,�<B"��.N$��ng��2tw0��$��}<XH��Rg3��,��U׋�!HmF��r#����RN[Tlw��R��
��x�TT����Q�68���*,��eBg;5�r�=u�&�uW�"Z�fl���oB�.�r�-�}1&Gx�p5s-���0��'�e$�[�B�4�ً(	_�⋍�_�"�v���f��Ge��ZS�F=�N�x<j��A s<s���+��T����H�.���Fj[�=#k7��6�z��R_/��Z�?*OxԳ�"VCRE�eH�1w���?���4�=��D�h@�T��k����&M&zw���V�Z>���q�Ϳ�S�>H�4A��t�y/�A�;��iNG�h���Wҧ��[�b=�.�S�@Ӈ���J�;A �#����.�Ugi�Mf��h:��i�S�ajK�Ř�0-�B���K�.���Ob��B�7L!lp���aݭ�=2�(�k��mn�+	 �.[(���dW��2Wb?��%�U9޹Q��S���ƘȀ�v�%J�0}��C�U��i֓�U%��x9�T�`'��̉:Z�2*��,e�`'z0���\��(?���HA�6�(���0��?��n��/����O����Ŝk\�X��Q�KMn����:��%�ɕXGe��f�����,ȓ�Т=�����ò\��:�ozqA1<��	�Yb)�� ��+����9�og!��g�x�8���d�ŹL ��B�C�TD�1�ډ�(���i���> ��ъ�[�e�o�E�8����S�D��й�7:�I�{����ы�J�E\�ؤ:fW��-1`��;�,<��o��Ak%r��-�4�0"��vv{�k~A0�����h�
�꿺�~�{�! }�+���-:�x�)��ڀ�粿G����@�
�@^��y+,�w@��O n��`)��ʯ�������K��=�UMG����̮L�ߌK�rޚ~�>�e�i6��Z.� R����i��	8(����4τQ���$B�"���43����k�|�!	%�Or��N��ߖɗ��;��D%w���|��3-��� ��n1�d#}�KW�@P��� ��*��)�r��1�$Iʼ3�뀮�S/D.L�(ǘ��B���{vu<��h�u?�m�$y3t��h��7C�R?�[DE��ԋ\�d�O���l���iI����5��_�I(j��AU���X��8��*�O� �>�;�f`<{���4m���Y�s/��4�_��cXw��H����h0?A�AWH���U!CW����L�\ɻz�Z	<#Ol�nhq�C펇��.��8>��A��
_�4xX*�Uݹ2�ḙ@����� �4���k��L*n����9� ���צ�{N��n��5��!���'����;;�*��Gu�$�E����~�}�-�p�;���?�}&ul��6<����	�[���}����^��CZy�t��X��Z����
��8$kS�`^P������ݔf�ԛ!�3��6�'�A��ʰ�
���]�Eɿ����:�ۭ~�fz<s���|��H�Ns�UCb�lM{\�7תBD#	�;��/;WEpb�k"����0خ���np��Y�6���6lE�z/o�V�'�	��y����.=:�͊�� $�'�y�Z�h�.9�8J�f��@�Q�:������`k�ctwS�Z7���.3�ď��"Ƚ�}��	3 m�����j��s�����	@�|E3;�W,�����D�H���2B\p4��9:�4p��ñ�28s� N_H��8�������"6��۩��U��^^��w��y6D���T�4�H������w����
l#a���9g%�t���a���=b�x�̅3	��^0؇��\��6Q�n�X+�{'���TȜ�lm9�X<H ��kȚ���eKd�R0�C��:O����ةx�$�W�7�N!�;��c�f�
��@V��Ia��`6�D��t��3����F��ۃ]KJgQ�q�粬�d_�9" µ�n"�(r�v����zs�'ڗ��'|b�1��������ӈ@��zK'hR�E��2} ������y'vX�c(Y���	9P���*���_��-('B�<Q)'�9H��{��"S\N�[J�e#X� ���{'q��?m�0ʑ휳q�б�?	č�
bn�� �^�m)k�1`�*���-i�rɄ�
���=�t�՘�.E}֔誩�&e���r`��ݵmFi�pїuG�AnN2p�0����Q-5w���~��t�A|��>_A#�
%0'����M�ߵ2�slZ���rK�Kn�E���	��{�Ma���y�����Tzx�¶$?� U�W�F$��m-d�'4+���B|�2ۊC�Kc-0|e���Ӑٙ~�^��@�w^��J�!H�
82�jAǅͯ�&�	�y�A��H�T�ά-x�;`��)�b�Ɏ�'���YP=Y���Rn���g��� F��C�B�݆��K_N��%	]XX�\�,������W�w�5h���m�$���߁����i<�`�M4>�,iU�A*38a�5d0�⏓pr�/��%3f����\���F�H$꒥��r�����k��к�u��Ct!���8?���g.�`�2�j���ލHt~x�E8����L�C���ao�
�N&L!@N��y�&u���F�Љ�L<��2�0�s�o�l��ޒ��Z��xJ�6ɁyN�X���(G����	�m��I�k�I��zq�?H��g�퀾�H��vI5�~�+=�X�4��I�$��h��8F+�O�7��ӻ�@R6��ّ#�a��*�UM4��Pj��X����w�expi���N��S
®J������ݑ��
Z��$�|+H��8��1��K4oQ*��{0�U����Gf�0���,�m��3�r�躯5�Z�Q���)iӯ&�� ����t�t^�Ӥ]�AyQ��(�E~<dQm��Q!!.y�[*UBh��j�;����i�r��B�����GPz��EF�R�
jj��nw!d�MM��^%(Ii�4BI6�W*��)��T�[;0����oJ�������Ԙ�&P�]*� } �5�2Bj���3��ҵ���b�͛�=��=��J1ad	�v�³��ؕ���T�:�)��-�x�TV�Jb��E(�J��	�ߒ/��HnT��[��8p{�Ux�o���s�ϟ5"�j�r���V'��p-ՙ]�/x�Q�.�7X:2'����^��?j�/��\<�~B�A[�U��a+ 3]���F`��6AN�_�D�]��-s?NA�KX��3v֞wYqM����i�;����R*٭#B����q]B�]юtn��%���oo���l���e�����nfI�R��Şj�#mv�ˮ9��8:��1��T�G�1������C�1��P����ή���=5~^��@~Z����ɿ͢u�L�sov�-��h�J8�s�p�b2�l�Q�ü{0Qo�i��R4��H@�xV�Ԋ>-h�3��2����l��.X�f<6ŚR������ ��;��&�ZL�d�����2}V���~�������60g�z� 
�ď��e5��3�02��0�����E9IA�M �GfR;F3w9�b���G�(@�	� @b��2u��r�d٠ٗe�/��������u�9!�J⃳M)<�����!:XQ_,�Őh����1��Z�t@�;a�e]��C� ��������U\�GQbG���0�J��J����ׯ�����}< �(ߣ��O�������92H�g�^42��}�{sV���+i�E�����Jo���@B׉"�?ضV��H�������7~�S� ��$" z����^~�ⴣ���Fñ(p�(t�����҆� �G���6����.������ȡ*vn�+����/5)
Z��ٛ�e����x�|�{���m�$�� n�i��(Ѳ�=K!��n@�����	�`�!Rhl$��?����T�2�O����Ou�c�jq�m�c%�l�6a���.L�X{�fY^gw��0���+������;����p7?�����x�܋eh�ZB�������hDt6z�8�A��8Ĩ��{BٍR9�̎��U�Ǚ��Y����Iv|\u]����wK��r?���졲=���R��4L���&~�uCw��4���^4:������o3XE�< ���ԝ�Z���4_eVPmQ�M3��w�G�Qݥ�Wy1�NQvs�L�VB	�Σ��C���Ć�̬�^������ڗ�w8Ł��`�En�y�2r*[�w���U�w�e�4��>v�������?M����V/H���n��������iL3|T�W[47���މp�҈X�k�o�f���:H�
��F�>�#"t�����/?���4�}�{E�}׋":�${����H7&�O�mK��]�|��ZW���h3��W�H�м�E �.+8����i}��Q7�j�S�֟�*(�ĺ���I���z3����m@c�!Bj�+Oªa!;�9Dj����R���f;����=c�`-,F�y2=������hh2�Kэ;�7�@�~�X�L7�H�t�����2����C3-�i:�K��\q�j�;�zJF�+��WJ%�@�x[��Ć8������~Lܽ�&�ݬ��cԃ$��5ev�ޯ�q<�<hm��c{0�^ǂÎ���gzq�,��?�R<���k2���r+���v�B���U����ψ�a�vhh���"i��+��Z�t]��������N3_��t�;&Ν��V��N9)+TP����~3hQ�~ؔ�!﫩tb�u�g��C��!���� �)�.��rt���3���9)�%���g�cb�s�A1�������Յ��ܴO�pl��{T��P/��mBB̉�_��=G̿�@�L[q�!��L:��p70l�T�%c�XO�	jF��مH��r�8cOya/�W2��=�)2�^����^Vd�� ���S�J�����T<]��@�ix�"�y����L�L%~˻��-�0��5�œ��G�wp����9�*�$A'������������n{
\��������B���8�j���G�c��}����dW���PG��DG���$���5�*�w��Bf胊�ȕp���u�nR��6W� �~�'}��3�Z��#0Ӵw˧�N�Kcx�CY�Y�1r�n�|E�'��h"�lа�TT��S����4����ed���xH�\{W���t�ӰO�ۯ)�l��@B'}�H�3yj�T��IK��l�I��ʲ&���Җ�o���ԼU��C�36��Aqo�s��50ʞ�?�..&ν=� _xD���$��v[s"C�⠒".�����M� �-�G�/�kL�DE�8��wx�CF��w#W�NZ����3(�+�<o��ٌ�������w�ۀ�MJ	u=��b#�?���ZI�`,
y�Ba�xŁ��Eg$��m�wDi�3���Ch�E�qe��oD�(�hV����2rܲ鏵���.�]I5tLH�}5��Bޜ�zj+�w��	!����%��*P� 3����~�N����F�(Up.��nݡSWJ��>j�`�akG����B�I�*!t�����l�P�M��T�!@RYT`g��z�7�-�\�2Ȇ�����k��ɩ�,G��F�LW{/��s��M ��jy:ݗY]??;Z�N-qW׶�!�������7�pd�3ſw&���uHZ�_5��,��Vye��OWB��7a(�l��'S�v.��C�?�Zs2��sl�*ߺ$:��q�"� ����Zw�䯔�8מX��c�`-'j�{j�`O�J"nf�1��X���0n#��|�s��=
C.~ބ-.���v���y���3@L�Z8�H�^�!����Hٻ]��0�!�G���ԫz����B��X4V���T�y��?j��=����=:��-&t!	e,��2�U5�@N~u��c��S�:�J�Z�8ك�]����L�>kY������4�6����A��.������8��=!�������n
���֮��!_!�I�q�p�4/�I�]��C+��ե&F%��{V�)��gu��+�6��3���VgYP��*��W$��Pm���,�X�x�tCڐFz���� 0.F��'HܮZk�����'2�R�y��ܾL��ċy��-�E��$�X�#6����p�τQ��6�a�f@�E�{����Y+�]����j�Է:�x�/�`/u9��;�ܗ��P�Ƽ���֐<݆}�hQb�g�j4��ZūW0ܯD�y#�vTЙ�\�$��#��G���(�u��P��A�y��G�i![�o]/��T��e�9�_�1\���x>�'�։�<s�'��Ӭ�A�[������Ƀր�����z�y5:����!h�6���?���wZ�+����l�b���?s�K�����Mk�HɱIڤ�m:TlxZ�hc��wio��JQ�\/�o�=����@裎�2��3��D����'E��<5�	A�F\���1��S��k��(��ނ�zyTK����������X�Q؇��YУpc� �R�5���d�.![+���θ�`�i���}#uѠ�BM���mSri=�>�iݕI�r"��R�ReP�A��:�l���k�,�R_�S��h�;��C����Oؚ��u��<KP��k��֭:bu(๥E_N�{~ܺ4���M�;�P��P 22��&z�g�$a�!5O2�a��)��8�`��a����RH�Sa�g��<p"��m�ࠃ��I��BW3p~{��*l[@o}���)z���;'ų
n��=)�n��d���݋������T9������/�(xYV�{��(4�`�%��~����vcU_*ᴱ�^�1��˚�X���9(���Y�Ѳ-����r}���`d���;�Ca��z`	Œ�Μ��_���ǴA����4s��5s ��`�/���Iʋy�+ి�m�rv���%����E0/6ԁg�yE�N�mo�4�U��P9)��)�i�#�b���+��2�!��[FT r�~�=�;�����ҫ��;:����e�x�� ��о�w�]���I_��(j&�<���+?�yO�����P=kpļ�0��V��qf�]�vw����$�$�}r���O��C���_�xov��4�1����_�"+l"oA�f�8@��
��6��;������훶\�P�3�a���/��:I]�٘�e~'�=�L�̂˶f��<Ss*O!��A�I��ϒ������Q�
L���a��V���`��{�����2���G)�Y�#�8dSg�R�����(�GٶRB�%�U褞?{^����҉���F�6�� v6�$�*�7��NF��j�!��d�5?ܔ
���IU1�A�*��w��Ú����"��P�^�Ynoi��Wa�t�*�Ƿݬ$i(#,jH\ʵ���'�Wkx������5G	^	!���:	t9����I��T^Jb'���*��e1�V�+�D�M��asx0���g8M�S�iĊ4./JV�C��Gu/�*T�iJ�WxԼ�M�q���I�v��CN����hr��0���xd`V6پ�MY��¬�d�e�Y忦�9��B�6�F��~��~����$C#q�1����|X Ketu�ͺt������٪�ȗh�b�լ{~ƭ��b67~�D��%j�C�vQ�1�4S��,i�p�3�<�w��<�8�c�_$X�=�J:��J�L<�vj����I�fa���A2��=�0���Y�w�=��Թ�~�� h=�Pnc)�ǳK�r�c�$ڔaE��uT$Us����B*`���1�8��#t�\�T�\�E0<v��fOPk(��fDT2V��p���a��xl>a)L������;])���r�%L�L��|�� =/����VRT}՞�[��B�04׿͑�+/�؎ɩ>��ϰ��\Ú��z��c3yID�7������YW@ߚ+��ѼY���!��x�F�7�z���[5F��6`7����|h�f��8����k>����*�.��>G3�9mo�#��yĳ��I2�&�Pu �@�s��e��j8X����-��!<Y���er>b��5�k�9�%8�P����E7f_9�[�qź�tּ�pP�����-�q����u���``z�Q(ţP���i��>܍��X���:��T��]#̰���$;�*9S�b�8����j����㟍�2N��H��:E����3�#����B��l�Jps�@Ǔ��~f�ǆ���3�$Q�U���,�d����R��dzk�O]��:b^"�=�M�*��'!:�����t	�w�:�Xx�G��`���m&+���A�*�Ω�?S��mҫ@�X��z��w[S�>�q��	���#��ZP��p��6̋`��n����3�q&b�	���F{�Q� �>&06<�{�MSG�.W0��5oe��DUA�If$l3�n�p���Y�]-�yҕxN��Ͳ�@�6qY>q��ѧ
�R�&�#p��ˬC��s��F�r����j��S�8�f"hi������o���Lќ��ؿ,��7��A%�����{�$X���ͫ=BHZv.�$]�_�&�r�'�� �������L:���6�
���|�vp�k��a�ʃ�w���vXq��͘��2��>��CR7?��?���)��qzYL0�����*���$�������K�LoCV�K����z�Q#A=sQ�K�@,M��Hp����h��4��ܨ<��`e�d�^v��X\9{2�dCwXuwT8�����)y6'��(������Q�SL�R�o�Ν�o9�ړ � �/�¢��C�}n�	��A����A��f�J�us���N2�D�58����$Z$��.�ٸ2q���>3��ۥxT��Yy���{�W��	S�ŊG�{&�g����=�d��
K�t�$PW���η+S��09�˹P��V+���G��x��@3?XW�\�ϣ���7��O������[g(����o��J*@��"3�a���&�n#?�na��r����	��H� J�U�a�rD<w�Bf�X�[Gq�8n�[|ЪV�S�6��ȏ�@`3۫�Bg�52�Kn]C`��̰�\�r=U��O!;��}�|�\5�C�J�GW $�$ǯ?��-o�� �v2
d�o�Z�<�@�<΅�A˳�j�vE�l�(�t�|������j���~�7�ϓUcQs�K�E���]�	&A!��zE�dUO��J�G���Ԋ��*�p��P�]���`�*V�p�1]G?���R��N� �mb���v��y��h+�k?�n���	7��e�v�^�$���.1�w�pF�o!��QM����~PJJ����;�,���a/��H�&��V������}V���*q��wp�X�O���>c���b�/���|(l�)΁I #Z��h�*�Fn/D���nPH����%�c]N�=.��k7�
�����h]�d'�J���s��8RkI�?���=R����ś��B�i��\^^z\�~ɾ�1kD��lF�l}F-ia��x�\r��5Tϱ��TZ������5c��P��C��̍��U�i�D3�5����:�o��y����ϒ5�UE������l���?�>��� ��"����}��5�n�� c�#UZ�"w�)4�K3�M�M�W|�����x��쑚fk6	�*�[��;������BV8�}{�Ю��u�j9����FKV��4|�+�M��� .n�}���^r �6��U�V�����~N��]�l���|�oc�_72a����W����CS�B_x�U,����%R͜f�����O��Ў�g͎O�۲n�e�B�=�/zfw������((!�Df�Y�X��Y�c�b��8*O7 :�<�=D	UÊh��0���0��
tA6$j�]$�#U0�!L�[RS�.q	�� �� �D^A�p��KU8�`-AU����UD��סݵ��=���E�ђ/!���#��eW����������#4�<G�K�aV�]p�9r��%tXe��*��I���F3v���)^�RH+�,����U�Ρ/�E��94��u�t��ĕ��C��N/h��s�8؛[�ħe��:�b�?�I�����ўX{��܂x1Â�qub����'����'�Ҍ�Z

_��^M��"�}/�	80f�d�f;�!�V�j�'":j�M�5�ʂ)L�T�:�s��T�Й�x���V�࢜�X�|th��Y'O�B� q���f�J	D@`�t����z'�D���[L����*����?����բd	�.=>7�f*���A���_|J����#{)V���N�cQi�:�l;29�[�&�F�UL���t��n��w��DX�؎�r�N�2R "m+����ډ�Y�W�F{�3b�z�e4a���%���)��������zO���9���A}��V�-�����>uK�
Q'��w�n�e�Hu�Ɔ0;�8�≥떛��mr3K�;����N��ލ���k�@��e�e�T8W���E%��[%�HI+Gg��P
�7(k�rf��h.�I�L�=,���ἿoB����ۯ�0tykdҳ�}9 �~'��ė�+D���I'��~#����������l�cZ`�늽l��"}�R�
�\�E(	�),t��y�B�����03!1�+c�Q19�1Rj����0I�e,7�y��cI�%5o#����kV���񣅣�|<@W��Gj�]��R�wu�Aܙ��\lw��Z�si�CBU�٨���'�%�#h=�r� ��hGO��%�N5O�X�N)W<6����4w�S�ic�y]�vCYtV�+�6_�«�y�	y)��-H��MX��q�y�NJ������ȡB�ￛi���4�*��1<̟���j`>� 0���u�sw,7}gIc��:���Ql�9#�B������*\�M����ŉFbi��A.����ġ�D�[�\�\��h�����t���=S�״�]���)���:u���$$��U�7��;�Û(+@?�-��N��A��|�>���S��D�{C�W�?���_���Q��,�t���q��/���/ZN{��۾�@K��͆R>�
��<	�²��J�вB+pZ�x��*�8?ڍysb�� |��M�~��j�6�����o@NSW�������/�ԃhP a��4`��/LG"1�jO�ya��/j!'2e�$)]?P�+��7o��+�����#&W֝���|G����8H�J�*�0C��f{���N����i�V�p�I7�"K���Tᝋ��D\*0�vؖk\ ��`	�U���|N)Z'�?�Hqu�d��~����,�#��B_� ��I�97`��5ʜ�	�L�u�hlg]^�2Ԍ�Ck2�1lg
��9�a��#��#bH���E��Px�x�ۧ#��5��_�+���C�^D���WIL��/.m-�j8��q������s���8��M��pi;�̓.�"Tf��4��� x�L��5�#���_W{�bG���W֢E�����Y�<ܝ�RW��0-DŖ-ͻ�������oܯ$Y%�7�"J$�ʹZ曆��D#A�w���w{�DTŴ�/׏:ԋ^n'譻jITA����*d���'��EK��wo7	)zf����Փ�D�OϬB��A�P���B��׾�MȰ�R@��D�zr�w�R��8�F�Ha���~\j�h�|xx��������
@��zM�`�y""�%�W�%P�[[��Q��h���~)�;�H���+H��P����PMl<�\U�"��J��3L�6"P��=)-�Wg��-&z_n>��0	��7��R��?�P��s���SX@�v��b<Į^�N\��������g>�-\�ȳ��%�}�fg�����S�����0yl}.2ǆ�����YT�"�ն,F��r�	U�"f����9Qq]S����4�[��@)�� �0�i��<�7�e�t\�k	��}�hd��IB�F��$ϵ��M-3�o�Q,�r�;qn �1J��Q���-$���jV�4$�yU�$������⒒��䉴�j-<����O���܉��:3U��I��G��o�P{�B����`M[º�qW������h_θ�\o������"ߙ��R�2�޲v�%�1LȤ˪Y���4u�W-�օ%�_��T�^\�����!�-*/�rI\�7�Ta�r���;�Cۘ&�u��S�~.ȝ���O�ԣh�Y�T����Y�=��c��
��u���g)Cb��|��5���_v�s���M���W`B��d)�57���x��/�@_q�� ��uD8�H�k�J��>'�!=�C�g����֧��2m{�"�G��?J�l:��C�F���:� �m������܅uǚ`)���ގ;��I0 ��o��n6����q�g��4�y:j`tbZtB�q�V�Z��V�����R������ĺ��x҄�T�"������@CϨF��s>W. Cʸ�lm�u+�F�>�U�ಚ�d�F�R5% ���Rd�� ����>~��f�cPg�B$V�$7��f6+�Ϩo����#v �N��8aeq��z��15FЅ���?�#I���|���
�](����i�ٰ��ҡ�XI��k�{Q��T6�~��=7�,u���}�I�Ĵ�U�q�����{o�[�.01����j��t��թNlc)�r�P.��+��]\�^�3֎;/�.�Rd�
_���-�;���LĚ:�^�����^ιp��� �QfM�<�=_"&�E�D
�A�;{�f����H�%?"��^W����k�Wv�c����;�MA��2�J,�����ͯ����z��x&^<ё�-���X� ����DÞ�����H�C�v(��|w9��)�M59g!��'S>\	i^�Gn��t,ꯉ��t*񸧊�8��x)4��!�"k^��s.N]
`�v@�� �?+��כ���J��R�"�a����n�g	t�I�aJ���<B�zSʐ=>�H���/�d��S��uёŘ|��E�AK/KCK*{]JX��*L�6G�<�4����;`cy6_�MP]Ʃg����g��!��埧��mb\'Gw���9)��i����G��� n�XQ���bfA�,,�J��T��`�����)�'� �{iq�D�}��@�1���k�0�BP�?�>!_	�nM�3͗�)��%O�v����o~������(S`X�HZ+4Ҳ!����E��u&�Q-`@�^p�s�5�U���Yh���^r}�Xpr� �������۾��G�q�E��I��aY�K��Ή��S0��Y��0�	����\�#�Q*�d�.?�����Ͽ���|
�ҕ�<�o�����Oz�'�'���2	( A�g�9F#8)�}|]�6;����#7����x���i�=d�jֱ���J��t����@&��Ɋ՜Y��nL��FW���	�b��`�t<3�������QQkg���U��*�8��v�������jF��>p[�L"Owzq�;�	IHyu�������-�Gk���;QIy^h>f�~k�& �|V�Q�����rp��c�깩~��M!l\і�.l �"k�����+�����(�hA�B��'x4`���E�*�N�u�aޡ��PY�݁�\A#"0D�<jgώ=�v%��7=qPr��:"��l�M���K�f>IAR�6�Z��s�p)�v��b?�O�{O+��_hn�H�Q^��]��+�eE_d�N�&l��:����W�h�ܯ=6�6��.��p�^4��f�^x*��_;U˿)��k�C�K��!��� U��s;^K[�v ���e�f!orG$���\�>)�(�ŧ|ޞ0�Q�@�|��sn�O�lY���eO�]��)x�f�&�7�؜AP�r�|�UO���y8H��ËT���y&7�*ͫIz�K�e�h)��9&�P[�.'�X���zK���,j�cAW/F�m���*� ��G0���_Sf�� ��q�c=|q� I�df�� ���Z��w/�ü覂�
�L�_!Z��G��@RdkIp�"ZoO*ͩ]�@(�X�����_���^��������b��"(x��d��|+�v�q�o�-X
q��{:�(�A<����TQ	�0���Ykq4`�qci���D��U#�柍��6s�>��N�PsZ�2U�/&b�1-V6�o���7��xf,�0�p~���R � ��ӼքFo�zǸ�3W\�TJ��.P,�w��H���rq��޸����k�I�����o:�r��meoQnJ�c"eŖ^�ťf	����O�w��v�7��έ�ZZ\Rs�F6X�'S �����<�蹫�h�" 0§	���*MO r� <f�%?61Q���ޅ�*�5�9&���gy�k����6�ܯ���c�M��Ƣ���Ɖ� ��g��Z�:��iFN���/��T�xr��v�:'S.AS�dȕP�WZ�̿�|�K��ڥ(��AÒ��jϢ͢�r�%��+ ���~;A��d��� �< �vWYi���{��4����]�U�(����8�`��<�ި<�c�%c&�	�N��}��*�pR�"]D���_�H�G���LI��zL7�43~�ދgY���2�
t|�2�MX��M�ɂ�n�q!��������a����a��~�R�W '����d��c+��}��ק�I	���c�߯z�|ue��-q�W��T;1H�d�}+����9`{�+촏�c!�����3���_X�(�c������Rv'^��ۊp�+K!pJ��t⹬5�e��7T(�	r�xk	xxVPlw'�|�	���u�
o��b�0�ћLW���K��B\
��G����o��s^ha�M͍q�ĥYZe���1��S�'��'��,h��-�޴õK����a��Dp�	������Cq�TG��2`�.����
z��\�\]�ؾ�TgI���[pT@:�ƹ_��-��O�^�R!�7�(E{Ryʈ�Rm[>h��J���D�����^�LsD��#��J��,��0$��ש���46�n�:�-7l�X�B�?)���L�oH����:,�����J���<!�ץ }0���N��� �a��	��4�p�3qe���xF�V��Š΃{Ah��o��r͈QQcFEH�-7��s���`y���J���i�A���J2f]�o����F�#W8��U�+
e��ܟw�@�ԎY�pI,(�q5�cG'�/��2�(ب!����ֈ�u�����TC����2A\��1g8?�6�9(u�glF����]�����׷I�6�m�Gl'�d��Z��a果�[��S���E�Ł6�_4��O����tz����c�)5������h�>��5n�߾��k�6OIQՊ_����+�����q�A/t�8��	��1�l@�¡�4&��ޮ]�RhD4�!�y�w.�KN/�ɠ�W��{�0���"ٰ����!�2��^������َJP4x2_r{�F��^�����	��i2�L��<Hgc���;�]�QDG���u�3:w r|��h�l�T�汬C h~���'�V:2�cHI�"Ro��pX
���DP���y�����e��bATt1�2���H�8�j�
R��FD�H��rd~���H�Q�����d��ɤ{�yX�`�u���tJ9���8ܗ������oXW�~u����6�@��(�V���B��f5���{�zo<���x1h��G��@�jq��v�$��ƨ�y�.�	,�xz"�����nc���:�"%��H������K��4��暤6��Y!����@�v���^�K!�B,��YHS�Ot�K!���Rj�×s"�HS��wV�C!�h� ���άXCr��6�fη^}�ջ��|~ϹD��w>l�@CS��D�ּQ��Ԣ���>ʎ~��ȥ�8V7s�2ڭ$Ҩ����Km�1�����N&w'!̄��ӝ`��]�K��wE=Zz:$�hv���%�֋G{��n{����*�����8x�����2g����ot�������7���;~�2���؅��K#N�j��3�+T�-cET&���&����Q��7��s�n�Je�;�E�]Q<�6 �Z��Q|�z�UK�0�����a�R������82R�赕$�L?��JF��J����[�?��,&D =����/4dor���U��?��we�7�YY>�S�C��w�P�33e�[*,я�����?le�g�_Z�v����i�~�|1>H�t!��V���틼
h��@$����(��W$���ͭ킿�@�A2#D�Z�5iL1���N���<u_>ws�TZ#T{Cs�	�UTl^���wWyA�l]�A�#Ε'���$"���&4-�J�2
�(���c]m݁������D1���7��E2Z�^X�u���AhkT�+�g��PJٻ ��*-�7'��rCUn��UB跚i�����Om�4����5��}�6���6�l������.������2�=x걸�����"e3z���oI��S�vQQj:Q��`9 ��xj������[z�n.���3�S��S[%�ƒz��
 �<�h���E��$n�.�˖F̄bwnJh�op]W>wn��K��<�o�2�em��(�D�0A�;p���6&@~%}G"���G%��N�b�
V�? ������z�G�$W.�����&�Q%����*�7J�/�Cu�6^�V���<�*�P�����kf"�
�>��BPEI����w��o�P\�1)��;j����v��<~4�"�g�#`�1��]�:�Lh{�;���3AV!*F�^[�l�:��xX\��$�_Q���{���~���j��J,���ۨ�Ƞ/LB;kT�`��ںޮ-�W6lX���޺��Ь=�c>؍%��@�s:M�À������m"��b�B����R����o��2����Yæ�~�,�!�Qֳv����b�en1�!ĕ���z��MQAV �y��7g���'����K�C\ݸ����V��ձ��J.4�'L�eZ
�i4�Or�*>^�1���3uϖ��I�V�g�҈O�f�=?��X����Ŗ�Iޝ�V|��\�|��q����� �8
��'�
g�!����� ��w�9jY��+�"�]P�٫�cOc�>+��z�����[z�b)=�:���nƖB����e{z��i��.{&�ɩV�a������lJ��6�S�s�����|�O�;��ǝ�=]�"��Z��|��yJ���`�5���'��j�����z<Ȍ����_�b@����a��=������n9�LU˿�S�(n�]��aa�fr�Z���|m��!D���˥�W��FgAnS0CM�`t>���8;z�����+[]���@�m,�Ca��P�J�4$�E���ɛM�òǁ$h�&6&��s|l k֬�wb����!�n!���<��/��YTf��!������_��@j�E� :����cA^g�J#=[F�ճ�����h�+��"�Mĸ���\�i ���z����-�4���d㸟�R�6��FҰ��C�:�Ͼ��|����H���.�����Hp�"���ڸ}<I�\@������1����3A���%F�&������H�	�@�V�YgL��|�����	u\���У�T��[��7��.ו☀�A��n��f?�}��Z~6�7��o�_k�E�o��H	���!C���9E�VQ(}{z����k��
�y��x]ܩ��|16It�Y hA�G3��'R��j>�7�-�,9��ZO����}�?�(��p���ù�h%��wGZ���{ �;1Z\'>�R&[ȊBP��
��Vo.P�'����ۖ��I��>�T�[z���"\�Ce|�4��%�yKrҏ�U�	I�����[�����ģꄒ��[C:�@��0�yTԇ�m�AHH~ <�-D6�6g���7�����^F_)j�@��4 ˸�8ے�&O\�7�I��;%�d&���g ��9��Mi��=k�`(I�LeFG����L*��J. �@]u������%�P�En��(�b��,�ڹn��2�ԭZ�i�Mw��{�r$��*=h/�ѸB�}�q����ZD8Ôf�ĩ��M��%��G����Zl�$.B�Y�bhܼ�k�ecaRQ�$�4&�J<>_NH%�֓;z�ӧ)Xr�6D3e�]z
f"l��v�Z~z]d��U��$(#A���r}�튅B�W����9�VzQ�+�UL!�K�\b(ʬט�!��iX��j���9����.��Iۥk�lp�5Vp,/n啠�-�[�>��3���x�R��6�p���~��u�Lڗ,~��_r����Nl�Ȓ4v�ao�h+��Ria����� 7��,ٚW�^4n9�Sq�����٫E9�Yx�!o/Fc�wDD,]�g_�Ŝ�--�3� ڰq�x�W|�7o���0�C(�W��'_+4��;a����4�����/i�b*>bc�aB��͈:�`�)1��!�1� ��{�k{�����sN�1Q^�j��^Ȍ��E�����K���W���m�i&}����K���Y��Wlu-%*�����RJ4��.��9ِK�ӶF�X��/������IF}jo�w�ӬY	��%k�̙9��P�Ĭ0�TW9tmW�����(��l�u����e�k������Y�9�Z
$8������I5̍��ů�X�F5����	9��/�q`0ӷ,��x3�\$cZ��F��[�c��4�*Ħ����շ$�+�
(b�ϑW�`���g�t��]d�K�1^������S�ކ�j7���K$*��	ލs��hǚ���A@SXR���g���j�3���o���Xa0|��@V����� |�R� �7yB�c
�F�_�ߢL�>�VR2�h��Wn�t`v��P�l#�u�p�Li���Zro�C�^�����]��Ѹy�\�~ߜz;���'w��~���8x}fݥ������yЇ���M~�S��Oa)L)�=�p[���jT�ɿ���R�]�ih1�Mg�z�y4hmo+�J'X�����%�S� t5s�h�~�=s�k���w�m�-M�:�׬���)S^��\BpM~��QL2���=%»��"u\�ǳX��Km�2,v%���V��n�d�6�!��吁̀��b��1f\f
�M��E e�]�F�e_"��ү�F��j���;l~�l�و>����2xų�ҡrwW$���`Et�����(	�҂h��&/C������?���R@F1���{�$�v�l/�FQ"���^�jv�zhV�}�W��T��T_�����^���8��J!=N�7r6�!a��L��.5Aί�HP�ybTs�+��SNtq�'>����ٗ��4w ��A˳�/$$��2���'ZՕ�Q���(�Z61�2e8���3yQR��A^+���of�Q`�'\H0�`vϠ��<)h�de�95���s�g��E�\]�Ȋl��D���'��p��|�Y"���A�!E|�u\�)�;��=���%:�A��D���tx�r���\m����S��r��T*��a�j����$�q&0c�au㿅$���Z�	Uh$�I���u-ٞ�	�hi �n��O�o��M��{/��ܻ�]q�P�K�H.c����15ʼ㎩B��f��RWp$:��$'#��6�no�'�����^n� �W����.
gS�`J�T(��w�"=]���e��?l�"�$��cY�\�b�t������>�u�@��r�c�ɑ�_m�kؓ����/�|�b��q�؛�����E�H�^epv��xĄ���Ѷ�6�g��]L�$M_�g�3���i���hF4����1�B҉�r�ѯI�2�������F��`�j�<=k����opt���X^E�Y���,� ���^�}���.�,lD�#b����&1��� #q4 8�I)� K����N?�Ҧ�!M��)����02	��fa�ŏ��O���'�&�a�"�bz�sr�^~?L���p��~�3����jY|�{�(�wnX=����A��ª�x�n�jo҆�{¥�{VGU�Ba��#�����\`L\�0��"�G���;�s��.�d
"z1ph�����)��1����k{Z�����叅�?�z@~����2�~�|���*���z]yPi\�x>����;�Ȳ�M��	�
�K�L����X�p${��@�,�^*J�j���\G[��S>U�xK���OLǤ��G8�E�@0���gN8p'X=�#�l۠����v6cUz�M#�nv���,9���_|�E
�l�<�<��L�����J���+
m��]��<�}�<C�:h�5�Ha�h_*ɡ��h�:�g�
�B:s|e��ΰG4�`�
;�kJs<Q���/O���U��c-�S��xd3��c|�F�w�?}����ϩ:��4�M}��~���C�k9a�=��˥3�2Kb&]�:�]�9�����xe��˿pq���ݱ�	���m\��wQ��0����(�U'��-�a��MVBag	��l�c5��� :yb��<oQ&m���E=,�P��U�*��w�('9��b͗0���8T-�U�ޕT&���[;�dB��� Rծ��)\�#�@XDq. ����P�z��e#g�iD��Ѹ��M�-�m�b��Tߪ��j=�m6�,����?6y��?�hs���;���1�~���Ϻ��}������Y�X����f�}�M��&Rf�aT��M|2'P2e�5~ �cH���<�[����a4����N�,^�Ļ�i��tG袬�t�ɊP�����+�aE�k5��s:N������+���KN��� s�.�_М���N�q�D ���H=�!	�~X.�� �QP�O�L?=Ԩ�)��cig����5��~�Σ�4�kH����Y�<AV,g9]�Hy{5�˸Vt�_XrRRj""����O�0�(;�t�	N����W�#bu
u/�'�~SgVI���ݢ��s���]�e���<�v0)�w�}Х��d�#ߧ
$*0��D�S��rnh�hN[�Y%�{�G�`o�����nc�c�D]-R:��a�I�Î�o�����Ca����Q�B��2 ��j�P ��gu)`���=�|u	�A�*hU.�xrH&s;�zP���*����9&
�U�V�0Uv��C$
��R�3L�䆁���~��_��u�Vm\�8�@�эQ�j��D�01x����wv����3�	���4�k0O�!g��Vm$��~����h�6�<�P��d4�Ou�k='s����אr�j����+���&?:8�����^uXء�;��rc�=�iֱqԿ"nKA��p$p%��̑��D8�\���ht��L�V���z	�l���Mڭ{Tgr�ɕE��c�����qi�İ`�٨�;����������S0�q��l5�)}���/"����N~��y��V�-/Wy���M��.��5o����1뜼�'��`o4渭�5E�)4��uxLS�(��N�EBR�U1��eIg�o"��uf�ٽ/��Ҿ���4��"2�ᝧ+3����-=Y��1��[�ő抴�_�?h��]�Tٰ��:=#�ϭu���U?��������\�ׯ\���{�4E{�����E����R-� ���3�c���
����}+�l�T�*�!s\��#Z	��u/��L�5�>z��ٔ��K�F����ve۶ՍK��-���2Un ����>�y!.պJ����Tz����&I�z�CZ�̄vsOq� ��{Up�f��^M����)�-�(��1r�A�͏d��{-��R�k&K �I�p�l}{-VRaM+���*��ԧ��{����j��M��Y����ς��2��4�?[8�$AV7q+�U�g#���g��0�1e�o�cc�����c���Ϥj�)�!ġ׸���t2�
�_h��`�i��O�}H]�`~M������޿�>s�$a�r��[�ѣj@����}aA�AZd�q�~����l��] th�pڌ�H�e���'3.�9g��Bcn���fs獇01'4��92���9Ģ�p��d��!��3 ��Cu�'�H"�C�a#�|������ZB�O\����Ncoƣ��z3���L@.���̢�v}�ǲ<sW5L֟��� xc�˟�z$�c�B5�Y��� ʣ���S��l�N���M&�K��봻�H��¸2������]�����Tw�>w�$�ݮ*)�l�ɀ)�8���-!��}�RaU��.x�v׀Vo�$���LV��t�9��a�d�:��d00��u�>��03L0�E�1������0�!�5�	�EJo����E��ll��;�ZIq�@&�'�)���"�T�9\���&���$����&%)T����o#āg;��ίj�'\���ײ�mc,�����:�҆�Is�e��4�RO߅#�!s_X
����T	3N���s�ẻ��s 5�{5��js���dm�p�ɷ�"�?��Ԍ+�L<8�����4N�yg6e��^�S�c��?x�y]Y�$8����7�_�'l#��	����<�J����}�a��B������,8���tf�����8�9R��� ��!;��]�!���әԋbr٢�Ùr������F������31�VEG����qPN���d�wA;��� �M�P�&ǢZGi)���%���dn/�<���ɻ�����É�>����>�Oʖ[�V>���@r!���`�BU2sJ	�%��xnH����D��&�u)eN�Y�l_7Y7������Q1��\}R�p��0�&���_W	?Ђ�@w�;�����Q���ea���m���%��m+��Hpe���'����FT=�-$��+�x�J�Ndt�_{#z��j�9y�I%gj=W��݆|�f���:,u���A80p��F��F�|���9��}k-ߐ�_/g�����Q���Up�a��E�̸Q���{XzG��#���iHE��}u�hi��0�F�a�3��M��zCS�֑��xᶰ(.��z�O�[A���C�f�8s�<�����z���8��P��x�lXw��9bc+��g�V=
C�^yj7�-�����+�!���VtOie�,]C̜�����ow�O��kM(J�	��lm����0)i����zV�<�
u7c\iF�L���9�@��8[w1�$	 @��C2�:���J�k3��U���H_<Ł[h��کg��.J���ҍ���F�CQ*���k�=�џ���|�_Ok)�jܔ�ߧ��oe��L?V\x�6!���u�C�7:onx=p���)�snhU���Α���)^1�8F�f5�IY�ɢ,O�	�9��%r<e��O�>�[I���#���|�������M�7�Œ	}Q��F,�9j�PV����C>��~���f���uY1ʞ6�T�Fp���8��؉��� %ǻ��o�`�V����������SL��i`�w]el�/z��tTN�sp�S����)��-�����KtV5��ye�?���Z�o���>� 9�3X�+q�[��i��:�.>�c!&u�^����Hu�
�lA�:�h�*�4��լ��IیnkI�c����Y���Q������.��^��>�ߩ+
Pf�c�'Y�1f���7�u����5L�1�d�Y�ζ�#�g�t��?�l��,e̣�L�[&3�����o�0��h�����2]���k�V�/��߷��cV�n��h�����T�
����*1C���R�1}�5�o� ��u<��Z��� ��aϩ��&KF�����ɾ��;���T���^�c�=�Vg@�������}��l��ȣY��+�7/ֹ>�/���K�y��=�t@\a�4n�d�MY<�X���tz�v'̤>uM�h�"�	�j���o�z�q&D�Ti���>x��*mF���?o_�,�B;�ի%���8�YO�YiV�	�Pa$��:�,�sBQ��៮Z�腌7�"SI(g�u#���'���s�:�%�M����ݽ�`ɝ��*�Q��~QV}����(T1��޼�\�Έk�l�m�%8��,-Цy�DM<[c�_�g,o�W��	�:��oq��f��`�|�����d�9��wS��F���AUQ��ߌl��-�vi/�L��W�6ǒ򖐉^F,gt��믂+j�
X��F��[�P�y�]��d�L�Miƭ�׻t�x��e�P�T9�zq�Wv
��Z�kZn���ih���S�E� JE��A&���	J��������%`�n�b�B:��U9��C-1�I6,V�CW�e�\�R�@�j:��Y�J�7e���r���dP��}��R�j��N��@�]�x~Bٝ�7��a��2�G��j����qO��g�C$g��G]�W�Kڝ���9x��5�.!;\��]Qο_4-�X�����eO�-
�`%N�~_&>��}l�Jˁ� ��@�\�tà�M7�OM+���@�Т&m4�w�� �~�ў�BI�Z��of*�,�4䇝�P�6=E��v��BRY[M%�~�J����A#g��~�.�\�E,�ܾ�d'��z�_ϧ�9l/\��S����F?�f�T� ��K䉯�"pX҈����&�cӵ��2D�h������>����|x���2R6:]`"��Q���⧅�*�<b��p�x�q�Σ�a7%ͦ�X�cܻ0ĵ@�tF�񗣛�����iꎽi���_N�Sh>�~�T�l���ʢ������p���
l9����"� �NVw5��0��<��Ƿ4��/���ʼRm�Zi�^
�t.������h�i��OE��,Fx�~%A.g�9�i�2�w8�hd^dP������
�C+F�$�j�]������K��u��J���<�T�دu�\�t�,㎔q��{�
w�'��&�:C]xt��� ���\��=�ڟf\{.ۗq��w;m��	Cp�RXR�J��:Ɠ.A��n���+>H�1�`'���v�Xji��+c����k�_:��a9a�Q���v��Zh��}�_��q{G٦ ȴ�w\E�*���A����ƥ�Ceޑ�#f��T� ����y�=�]���t�u���p*J�5�ED�[:���#�PʲR@��d1��=��D����㝙��Y�����t�ƨ�{ـ�~���}����Y�-��f�;~�6<�q=�{{u2I�ۤbm]�`b��U�#i�zK�jm_}jC�t�Zӷf�t$
U�L�a1q�$Uaװ&:�'���A,b����"��A��K��Wݘ�d��E����C����@0�u���(d��A�heH�)�?�sYM9�!O$���|qʒA���B鏃��`R,��0��8��k_B'L��.������ç��{�|H!��:��е0��v��q���~8�S�è?�iEm��زD��<�հ�[�ߋ/n<��7m�SHF֖��v��Eb���Ҕ�������h������s��G*ڟ���X�B?.w�q�r����M61+������y�\O��� vJ2;:��A�1[�C0��O�e�W ����_\����HE"O�Ş]ҼA)�!�a���(y9Ky/����Y5���M=+��~�oO:9�{���ڵ,yM��,9!{.&�O���p1ԆJ;Y�f��C���@[u̡f6.Q$a�4�X�2nw���Jn�3U�}puP\Ro���c��N_�lx�"ޡ�=��f�yX���G۠�"r=�"v��˜ w��A�g�C�L��a��5�oKhu��%�&�rt���*!�pTjٌ,jF_�Xe�3�i~�������Q.��`Qӛ���Y�#����#�U�Ǌ,ٓW�;�h�N�ab��S].7`�H��*@Z�e(ۋ_W��M���{"�S��N���N�f���jۈ����������[6˚�EO(!���).��*I<�k��Y�9=V��6��2y��Uc-]���c�'�O�d>��H�l��1j�����Zf�f�d���7�k6
i��^����@�l�ba�$,] z��u�d&���>�l-XVG��DKY͍X�L闼U����G;!O}�O��]L��_�XIHu�	����(i�e^�\f�L���_�V�s� ���<��d?uϡ�ޔ��k}���{��l���]z���cY�
5�͑�v��V�e�w�M#P�_%:gG��RM��l|.���$*8�Q�C�ł�j̺��Q�N�\G���i��-��e��s���f�$�#��ʬ��n�N�()� j�FT��V�7+��EՁ���wm�=�S�k
gQ!��k�s�A�������O���ü(�3U�-ջ�7�(�_4ns.|�Fi%��
t�w�n��" ��+�L�����n��ni�di�1�+b�Τ�iŒK3��oȓf�\�ω��r�6��"�䴐,��AA[��[4uRi+>����W��R�9�J�/�L��kڍ�(Q�f/�)^����R��z�ͫe�~���*X(;�Ko~�f˩��5���g��O��wҳt�� 5�U])�v ��b�T��w}��*�T���	r�D��|`��a&��)�`e�f�L�0����D��L.��7�0����!���mH1NbP�=�t<�A�gD.�S��'��#Ė�@a�� �8�WT!��;M�����{D&�k ��L����r�[�~{vX��'�tM]9U S>>��"���2�����`@��]��������\o:��*�[,_��:��{��u�N�mSP�I����NyY�U�]����Zu��|�g�j�� /|p�Z%�~�6BZ��G/B��}���`E���Ӻ���͚��0q}��g���,o�C��,��a�����ʛ���x�U>��,����?㴤��b�w�D��X�����R��t��<����L����"��:�R�+{>9#��Ў���H"�r�m���/Pe���!�X3k��} 1���lǓ��Y"~�@lac6k�+p��'�[[�?պ�
}���Q�s����A���B��Q���<p��Q�6���nn���,�{U��Kޕ?���� ؕ��: ��evi��wk1�}��-VH�0��� �BK���
)�b��6<P�"K������kTҞb���,N�0v5�;Γ�@A�!�%��t�,����rYSBj[I0�T�Yb�e�:x^���O�D�A��|y�V~��C�_Pzk`B�ϋ:P �B��*3�� ���,��t8G�ZK:���6�ng}�@�s���+[���@&4�� ����{8
�kIw��(×����<z�(\�W��mǚ>Ml!E����Hg�]�j���⛳�*���,�`X�t}+�Z 9��E��4�_�B�$����$ �|-��������6T2t�6�)Ƨ��/�ׅ�1U�?�粒'p���Nug 7���I��־Zt�m�9LÎ*�d-��mt��`�&\/k��
� L�Bs���ށ�X/>��~��ı�^+�Q�ax��#��������O�z�����`wht�&2��R�ጢ�������a�)��It�F�&|@��ȨU:��!����E�3�>Nh�G(���p3�C���[P�̗�g��{>����?�>�n9�z_I��8�_/\�)�\=�����A�/�u�|[$LS�l�����5}��D���Y�+�V2�*�|"�,��1BL -�6b4�������=�2ȋ�O'��n��ʀ�� ݈�Β*�ޒ�Q_�������Pd�gúl����
�!�z�Zna1ܼ�ZI�P����L��6��ٴ�kF&���nM�Ob�3:k)t���r�P���g�Z�L��v��8���aɩO�t���<��͢r9�%q�h!�%\������S`�N��dr�c5�	�l�k�-痼����-6V˃�Ϗ��\��(�ąNS _��^}I╽4��rx�S��d��^2�`v<SJ2GR���-u����xU<�l%>��P�pՓ�@�JrJ:E�:�F��mY7��e���(��%@O8J�a���h�2�l$�%��*�=�b�����z�	0��L!��)�
꧄G�S%g�n�e�gC���qp�����&�5���'��|C�-)�W�F �gM�3N�]��ԧ=�ȻAaX>���&��Ț�%W0�6^`������{�4)O[	G[��	��l�b�#Kx;��8�?.MjH�	`j�a}������j���[蚌���4C1U�}!D���+�8�b���A87�*�{ݖS.V�)YԤ�F��?�g��Ȋ�随D�.&c���f����x=���6>0����"xe�v�o�Nܺ�#�?�����5���� 	��r�{R�H��w�ϗ�ӂA3i��W�\̛r�V\�k�⬸���/��b�+\�x�4yXhd�o���uk�̘+�x����T^�cZ�c(��ㅻ��>��IX�
��"��Do����R�&����s9eE�ߝ�\#>i0W���0�n���Mm���>��2��� i���B9�?B�[���?�"��xN��)	3Ƀ�Z�YV����c|Q=�OL�PZ�<
D�A��#�Va{Jd�1i;�N�1�1��[�K��HR?&"�#�&����e��BY"�=&sLzii�$�|���X�����uP��J��x.s��q���ӻ!1��ǅ$`�S�XF�����w��c_,�]�8��#� �/�(4撶+���2>>v�'��7�j�S-DF��-���(����(�Gr�lJ�e�rI�܆�^�*��m&&�'��Q�*y�{$~X�+��o��[O���k�s��n7G�Lc�	�C�^M���c0��s
�}8�0F��:�B���wNokh�r�IZ�I�@Wb����ŰB���Ҡ�͝Q����~-��3���=�����߃BF�N��CŲ����T8uX��S�H�A��+?(`�X���.����,���+Un���;}�D����
"�i���3ܳ�+�!7�#���Jx����̠>
d[=�Jg��t��K{�w�� �jJ<���$����v.f��jc��y��w��P��E�P+�e��E�>�<�^Mi�/�RhGFҠ<�#�����D�V;z���}+r�^*�W�l!p?����I� ���Ґ���-��YGa�=��>oT-����&O]��l6��4�*'&>��ӅwP��-C�>���"�_��<pc�jOl����K�?g�;_�qR1!��G�^�7���B�aG2�S����<Bʳ�(��1QBu��r3��^�_^\)N��ٳ �{��룃���m�/��1Ǘi ��c.Sʵ ��n�MwZ���9"��7���B�^���a>)��hj�l-�	�\@*'{b����+�+-���9=x��PL�xp�M�ڛb��2: 뗛�֣{$1	o��Ð|�����PF6;�Qq~-�3~��&�ԃ��.�SByI�cN浲�����`�e���B���V[�c����%�|8Y��x��~��>�7+pY[��"�_��0����8�\'ހ�E�K�(�Q��t6x����Э+���N��~�0�WĶ����4�i�Z�k�B}�P��4�hvD&�&Lb5Mr�,]�˗����/��n?���*>(^4#k����C�P�4��Y�t�jye{�"��[�iy����§�ك�ܾ,�D�a���lql�eHr�W��P�e�>��؍&�éa�?��r?B�����P|�>5AK�OG��Ţ���������3J̗����I�6콢=�,JY7g�"��b;ő3毀J�>�%,T��0ړ���Z��&�Kl�����0#h#�r��*�`�g$��H�-��]�sE�^�u�����k$56��kȥ-���܂���{�=�8����I2YQY9:�F^�^9�͎Ƹ�k%^�Č۹߆�s�IY��;J�_KC�T���]9��U��Gd�
PGʻ��^�:��fpm����,y��%�O.x=��(~��ҿ�����"�R~��VN�
	
�&y�d4�L��Ph���	�:��Q�D� -�2"}Q��0�^�{���i����xB�  Ͱ����{�<�o{��\�K���]��qݼU^K�M����7H����ԭ���GQk=D�g_J�4�:����a��_^���.m,��ŐKӬ�.^N��S��Ku�� ����[L���V�,��ꃔH^0F����xZUd��
�d���I�X&��D�'�	���矪��ï�8l�T���{�2v����/�����O�;�g�Jה��8A<Fx�"����m&V��
!�W8�x41\��@i=�	M}z��7��8�y�v1�Hvt�W�g�?:�&���h3�@z1x�6��j��$)����7P��Gr�H����m
3�Ǎr ��q�.=����7b�X��d�P�R�ݸiN��*f-N�-�aH�P�DHH��)P��
����./�����7���=��8V�8[ �J��Q ۑ�G6�	8�p \�,�/JG5�����{+���
���K��W�4�C�[L!�?� ��A�/yS��#�O�Z�QԖ���cA�
i�+���Z�}��#\6BB�{����k(��I��q5\O:��β6�ժ��^�m�oړ��4�e3�í1+�֊�kՖdP����L�����%b��!+�T��ݏw� ����.UGc#�|)]u���q	9����K�?�� ePf6�l���rp2����ͽT��Q�YD�Hd�c���ot�&��_�H�
ߝe�AX'�����(�1�S� V_r�F�J��ё�D�TL(���H|֢ͅ�B��׃�l��;�6Bp�ˁ�7<�^n������o) �#�h�k��z���c<5Έ7i0ã�/�,��Z�\��;�����h����B��o�̿1��U߁X���D�ԥ�����e�\ ~��je���V|XV�3�Л��/�P��:S��D���G��.�!���,��$*��cZ�w	�&�ν�$�Y���MZg*`��:���̀gk�ĖT���q"�W�W�*$����5�t!��ȩ0vť7iӨ���q׻ �<���}���o�w��^�P�C�+�uq?[>��Ї
~[�m<�X����1���ކ M���\�EBi(�g���_Y�'-:�ʬ=�}�ې+F�  7�Pg�e��$�`��1CG���BI��AD1mrV��;�}#�r��8� #ծ&��������<�DQ�|����x̻���o5�F�L�#�SxOr���18/c$Ayt�
�mC�b�7豝_I�`?K���:h]�(%t6gɊ�!�R�T��� YI�k��M:�����L��얾Ak�:��N�q�js�Ӫ�'�L$�&b���X���bD����:��$i�qR1b�Bk|)|���hP�e(�*�:X>	���F�I/]���U��F���_v����}�� 8�b9r�t�;�#c_T�Νo���&׾Q/�L���'��n���&@��g�l���/$�h�Ѕ�=},K���w)�� ����j~mx��L���J�4t�hQEV�9�Q-��":�4:�-�{�^�cM�����"�-��7���a,�pޒw)h��H�
�����_d���Vu]R9��`��b�
�uz�i]�yQ����x{;l��Ć��rv2�����b������>��7^�Ȕg`�v�S��]�X6TH��o�k�8}t����3���ʆ�tY裂�TK'ڸ�g���\����}=�������S����{�8�Nc�9 cT����ȷ?_�x�rࣨ�4C�^{
"~$ۛ9�ףʹh���Z7ˣ�pJTizf�ߣIqJ�.�t��:����&��S�#�b1`-�,�{qX������6	�JaX�@�V���1���ri{F�tA����ĩ�Ӈz�O�0!@�#�R�(-��nh�j{3k([�fmV���t�=",���x�\f.�=�Õ 	�e���6,I����ˌ���	�d��d����i���gr�����}$��ؿ�K�>�h�`y:�?W��|�3���R�&-e�5��&&�K��;� d����fA���IJ�ht!=��_���7\�,y�����<+f��%����Xsuon؃z�Xw��mH����%~�oN��íh4`��.������lM���m,�m���IVcH���N�D��*���.�7��=��`�2�oZ��%�{`Jv��ЖT���3G�<_�o��9���W3�C�N�&Rr9�k8� ����Y+��EZ��Q� �H!���7k�C���q��E��k�iƨ��$�eֆUz��E��T��
�Sm괲���t�����i8�@���!�\oݳq;��Q�ZD�O�Xg�Zd��E��󃦨�k�+�w�t�9�\D����?.=]�"�\UI"N�6W�r9���Z=�<~�1F�{Q��]���)p�Y�̟��C�Վ��)��eY�'���@�l�|S�9m�߭���P�����|;��Pw��Q��⿻�Q�0)�,|�ww2�_:�v���Q��ph��l�:�8��X�$a��9���]G|aq���e�9�QI��{������r}m�x�k%�� �\���x ��YS_(�(�L��Q��NO���&U���Ĩ�w��o��	'�����7+�f��[b��_�;ʾ}��� )�=��l�@�!��k�cj��EA�������l�,���(S6܋�5:�C״��\�;Ȍ��w�����F��d��+��a�`P� ��L��K�7hK�h��G:��#;�׊й�=��6�U�Gx��A�e���	���}���|�	p,���/%�d)��L&�!�O���U�<r��M���"VMI��7O6�k�B�N3���������}�mL�[&��H��<���C�{�%�_%0�O��_�qQ��b\�&�o�����n�{d�-���Y�MAf��y�k^�A�� �B���B���Y�sg����dt�%�>�xt����� ��}b��M�HIo&CR�R��b��4�m9B8�wUv�;�u'�T �Yi5���y�LU������~y�,�+��W�����ߝ���l��X�]Tw+�0���Ϗ��.`;اz7&�ʹ5a�=6������C�ڷ�؄LxBX�(I�CMl�DLMy����$�(Fe%zcܒ�o�#���J��[T��GdB�}M~O��1�Ox��11c�y���W�~�c�b���C�4E7��2`V�CvV��RY�o"[|#f<�u�G$QP�);��Z#�%=�m�VCm�Zٳ�Q/J�߉ 	v|�NR ����~���N�њEq0�o�.N�kN����g5W6?�=+��lY!��'ݣ��07t�^�n7�����/�K��Jcp|�D5Cb9H��-|�@`B����]�p��l+kb�GY3x�Bk�n	�P9vU�c�i|�}�_�ЯAMR]�潈`�Kq�Œ ��9ـbYNYj?����e>Df�]�cDmXZ�q1��@dUb��q2�3j�!K�|�Xc�-�TP�����^�����R
�����Ҭ'����A{!��HsK������;�m6�Ʋ��V�
����f|᭿]�����D� ^Y�°���Ld�8��ɋ�%x�m�L�}�4eE,K�xx�Y���{�L�~"=�]k�Lp*�ˈ����1zN�ۻ�
p�&�Y�k$08:�Ў���]����p�O��/�+f��"htB�~o].�����3��-�?�k�g���������I����ط�dA�n�!y��C&�c>�9b�����R|ɧ�8��T58�8�O���e���a�)����DT���ʄ�'��V
�jL/I$}o��4�>:�9�^+Dn�}K}ǫtO�@�*X�7A�+9��6U<f|�
�N/2r)vvA׾�b���aԑ�G�hS�_ǫ�U�pѻ�����!�WOC�k�����u�Q#~=� ��<�e���@�=��Hf�N3>�U�]R�#�t��W�&��q�Պ<�K�6f¶�@F�as�n	���(�g�O6E�.��u�y���ޓ`PW$����ʒ��Wi��T�'5J2������+��� �&�ȩ��t̃�\Q�H�i����Ҫ���Ĭ�
����~�� �-���X�g�-�j��k����d�n�� �)v�:ͺ��4Z����Js|2p�2d�K���5� >#�P��t/�f�p�U�Y �n�#�� ʟQ6�޳�a��Ya��QUlu��yh��ln�߃J���A�t��D4$6ㅼ٠�Ĉ;
��uN�g�~�lw�*��^�*@pk|P�']b+{�`�Y�ܿ�Q}/�Vu�[!S7�Oevg�(�_v��/OG�a G���<���/P� :5���
��#���t�pt5�^��J��Y�|�K�6�YS4���e�>{�M3�߁#7�Z�S��A �B_V_���j?��ax�Z����q�!��)��@U���݊��㘕�(;?�{����;�q����q�⥮"��QPt>3z�r��USU3����O�@�FB��Ǉ��V-���PF�4+5�"�Bl_e�y�{35`�fO9��X��]�.b�0Fu�w��E!�)�X�܍{�r@d�d:뱢��H��[�ґ8�E��k|h�Ke���Ǿ<��@��`<�Z��L?� ]�����c���_;����PÈ�� ���G��ջ���]YҊqYz��"h����7{�ܶDze>9뇙�3� �q�Q��]��.���x���>0G��zF=�y[�����v|(���i��ڵ� ZOy~�y�1`�3�%�k�Ar��w	�[������6�������Q���̋,O�vp&ki��=�k�O]

 *����&�1�<7�kb��vd�}
o&�!r�P!��߃Ƽ�~/��(6=��sj���Â�3K�S��A�5"ĕ��S��u���)�oPQz��
{R�0U�p���v���cy�����d�W~�o��`����f�vS�^&#W��,���d��
�MD)���L���D�d:O{�n����'��y�5��Tj������__i���\+��y	��0����ϙI��h��n�Q�P�B�T�Vg�>��aF����7x%�
W�+���X�3��ƭ��*x�W�{/h�d�7*��MB�LK�:z��`����`�z�O�Ks��9�|��׭��?�p��F��XS���V]zO�_���f�e����!�[o��U��>��V�8~��-~����&q{*��d���
����i����ƍ'PH����`�F���A��_����uIL�#c`�~��q"*��I���S`��8�){2b��5�{�Ս���G��Ę�H����\^�r�����Z�i 2�Ϡ��Ώ�e�vMO� Y��>u�Bg��"��
�8?���t)��w�N���D���B�����;�!~U&��1N��Q:�"��p�]�ɠ��՘��	��p��"��/���-�\w�5��]�I�M�Z`|�����1��7Y��,b;�K�Ht%�ۀgPK�Kxjrc�NιV���0�9nG�E�y%��v�bo�>^�SĎ)ڪߤk>�&��p��̐�¬9���u�q}Y��#�e&[I�� ���0�6f��yex�t7��բ��W��*�~=�]�berVV��?�2�X\뚵�f��r�� %�PL����"a�JߚA������
���f\/���%x��[����ea&����?��b�����y$\���;gP��|��u�?$Er(��ׇ��u�~YT!)��JW����V�o )��=��	��ZnJU��S8\����F �w�0�U�M���m��6������wRB ��t=�_�>=�Ƽ�`텻�ڵ��A�$�p����5�X��Sd����}�\(XU���Mf�B�S\6p�� ����_u��d���t��f|O�B�$�"��?����t5�^Mb�J��i �z�׶���j$��@�CI�q¤(Z�q�6Gt
��]����/�폑�!������5z�$D�}-^� �Ћ�\��lϚ�����N�kRFO�R��ف����J}�A�X��
u_� �5������`�����Ë�PӼI��V�*Z�s�E['��z�,6�>a��Wl����ܙ��	#�GWmEw��_��]� �w�8R���
m^�P.?��)FGR�@��n�w%B�Ō�%8w���׏R�%[:e��\v��@�y�!5o�,o8���įm;r��C�9ߚ�e�V����`G�a5ϋ��c.uCYXG6��LM��H�4�� �6̋���B��mdFM�΋*- kN(�-��i��X���0��o�`�s����ᆁ��%X*���"b݄�Ye��v���Z���X�͖jqg�.�d�7pݡr��q���7|B�d���\L~�C��8)T�����#����xM_2N��J��eO���~�P\�B�l_ �;�D�~�@'��TS��5=��E�PdQ��J�Ѧ�)���6B�wn�>�]���8��W'Re�rg�4����%��[��D
i@,���w��O�T����*̡YN�^{�/��q�a�}�k�Xg]\��|x�0ÒZ�&��0�H�����>��+�]R�w�*��B���iN����j$��ó��T~��4 �рv���?TD�@��>�JJ�:� �	���i�|�~�$}뚐CT���l*'Pۢ�C-�=��Ey�KYϑkT(��{�v� �!~��[�/��O�*�wYmMS�Fn�U2��I$��=��0m��gf	��<���یs'����-�&׶öQzP*ߘJ���e�iץ����@Z,��^><�M�ݽ5�f����� BV�Lǽ�-V��B����&l���[�#�2��1w�:�mo�_x�œ|�V��|�e�/�㜝��6~@��7f�(��j�/�W���#�����(r����;@���k�c̼�_Ln� �x�0�>΃���y���a���=�{i�|�����i� Q0����}I�6j��&���@Č��0��x���~}X�2O����78>�}� �)9@:�x�����l%�K/�U^�=Z�s�a���/l5K����N|ځ��J�Ԟ�T���;X�!�n��4�捿E�+��u���X���z�㭒��H�C.�2W�x	W�pZ��ᷘ�`<��[P�@�\~ƞ��Rqn�dU �׼�l � (�;^ ���l�m��/D�>c����2c�>֫T��,�q6'�}fFd��*�	�y���{�����ݜ/�nd�ʠ�G/y��Q�j��E��{����9@@���C��OmY!�1q͡�@V6���ϛoP��4�[� }��5�Dq�;V�#��gSU�_���fq�>� w���$��8ƚ�6:�?1��ꂳJ��L�kr�d*�;�6���h���ae	-���n��Xy�'N���d!+�?z �W�	*�����$u;�|�j��C���X���n]��Ac!u6o�j�*NW�5�b�_m��V���)�� ��HR�m�:�Y�����T�Lr튲��/�q�@�nO�g��CB<o�`b���q��P��;F�|[�
@fF��ܟ��(D�W�����s���A'��M���mtP�n��z�%��K��c)<'����9S�V>���R�2�1�A���;��=��]j�a��6J�þ"����"u��B"��T�O�Vw���,���)�#{�Oix�ɴH�-�MkF_N�{�6�H��U|��wQBB��M
{�K�E�����r_z���|���v��-p��Sjf�=��ƽ��O�5J��"�]j;*+�����Ζ'�pP��I���з�-�Y�dW�W�obl��q�U�Z��:A�/�v��WY1��C`����J�fYMbY�GJ�*��T���2>6�i���Kʐ�P�<֛u��$�r_[�ϙC �+A:T�1�D�eLx��m��>�^�!۔����p��^�������=�#��t��v{��3]��T�H�����)��u�5p�/��>o��O�':4 ��M����/z��s���<�z�\247R����a��8M�t��@ȧ[e׹�jށ�D�d�|5�4��a?R���?[jB��ٴG諥��'����3�A`8����M�|DN������F C���E��},2J��"*�Vq�l�_���e`����U;皸��X�}�(���w�����(}G~�M����0�IB
7�uv/d��ڈ���g��_V	۱
�ok�6L0��h��Fy��8�yE��uX4o�!\��hB̔v'ǒ�ꏅ��!M��  ��<���7���ݱG���O/��I�����Z�(�:L����m):^�9������[��Bݵ��h�K�ؚt	}�I*ׅ~��K��=kdhQ	�s�>;�F��ۛ���)��F��64z�-��|%nҝO���JץEuj�R^���K�� C]�K29P�:�Jm���J�-{!'Yȼ�Z��y�Q"(.�����E�2$�X3�e�������|L>�qG��Jg1�n�]Uԥ������|傷3��K�`��D���+Oc04^x�Me[U=R+6�;56G�'��׀o�����G(�HX���fmO�]R(�@����DC;T�VΕ:���`V{s2�F�-�i��4t܆�8�g�Ui ��P�Ύ�dee��%�Z�Er��mpe�M�w�`l	?b�"���ߘdA�Wʅ+
���n���NSɖ?H����*�X�� ƛ޹��!o�#P�#ì�"K)F�
nyVXx1~��	�S��t�?U��/��������f�&\_l�YFG
Br��Q5q_�J�[��� D[I(3|��,7��8����f
4��/ֲ/�:y�9eە��eE��JO��O�&���B��q��E�Dx>c_����|hq��N�N���m��,\�I�i��ل�J��/ۓ�"{�R�RfKd�����)/5ie�ِl�ƙ�Q�L�T�.n��Ř��c2��?"�����+@���*j�0a�Z�\N�Lx�o�ݕA&%����fQ#�� }��4���������4�lZ��D��XF۷�).����p9qe ��|9/Y%S�+�޳Q��[�W��`����ZG���dj�f��R��ӝS V��]����M�3ƃ�� �O��J{�=���ma<�#5���r�w8~��I\u�h9�(ΑD��:4�vA^���kt4`^q�t�}&J��qʆ�q�:�D"��.ۃ�-ZS����k���%�6���uB�0�e����jDFr�dz2>ԇx���I,ѻX�J�tK���9���XD�h���n{����ʷxh����罊e�J,�ܮK�o�����,KY�31uΣe���Ʀ*���9��t:c��DY@5����_a4$�8&z��P�P�n[�S���y�����!b�V:H���"h�+���R�;ۃ�=|͟L���NZ+B*�}S�Tc�Oϙe*�Ol�	y�X.`]_����T#�IS�t/Ҩ��7x�lJ�oJ������V ��M|�$n��m��M��� �IXI>t����Lܟ��1��"�{1���P6�L�,�2��b� �U-qaNӳ8LV�c�Y ��9~����9�?�Q��^q�5�M����B7�e��vwJ����rg�J��iژv��%��9x���3 ��p�$��W�PK?J8��7���9cu��!�]FR���~���l�QQ�6!RO��%{E%u����1�(\D(���6]����fY��/n+���g�	C�k���XJ5��b굛�Z��G�@I�S5�6��l�j/�H������83�Qg[�d�*�|+9��^�	�؅�2
�k���I��$]�M�����WkxE=J�׵C1���G;i�3�
��d���|Y�sf��u)~�l��c0����꼻�%{U�/�ʮ�%�Al�s��47R�����p�7 ��9�ʎ~��'i�����Ӭ�S��W1�4F������8j.�i��h�18�!p�ǀ|��Ɖy��h�
Ć���(�@�S�^��
Od^�<����[����������G�$��Uɓ�3����\oˀ���~�Y�r��qG|�;�$h�����K�?R���3Ǵ�w�1	�2��{���(��Ԓ��O��@���1��j�
oP��.�c�e�F覣YP���h<��3�*��K�w0[f:���E�Q��3�X
Nܬ��I.+t"�@o~݃G��O�wѕ1�X��)�p�Z���+���=&��*~	_c����%���Y��6��`$v�Uw�\���~96�.�i�!C")G%Nq��� �} �-��-��^���,�2�$��Ƞk�Y�ni�~`ו��)cD�n�R��]o'���[���3Fų�Q���6;�-�l�%U�j#N׺߉��PϗMK��Sb��Ld;7�$}r��"���a 6J!�x��nr~����{q��X:3M]F�I�n!��m|đ�-��M5��)��łF�/uw�>�L�CP����̩�.��)i!�N�<$�~����!��H[h�<^\�س�}��ݜ��T�k%vWȻR�j��
m?0�������|,�q$��|a�a^����E�rZ�Lv���}O�H�|<�h��X�c
@�sR�m?��v�O# ː�U�h�N��KӖ��XI���p2��0C�w�c��W�v�ҙ��4D�P���,��|�D�'5��B�� ����� ��2jL<?1.����e0��2y-�c�lĲ?�+��
�ț�����9M�<�(�^ZM	ᄇ�%X��75g�C]�BH�H�i�x	��u����6�z��X�$o�.��᜼��t#ʞ3��^[�Y5��o�j�hD&�Kj�tK�r)�4*Ի�ąD(�)��S���֜��#{_vp_��e��D	�9��������fh��ȑ;�̬Ɉ����X]�2��lՊh(	zi:6�^T�%ԧ��O�#>��-�3������_?7:@q�|a�+L]O��)��>�O#��rė���c&�솳xdt:�`w+}�v�ܢ0jW�� ���;�aa{2�v�1��d�'�G	����#
.���k��3��#/_R-NN�>�4Nd�Gs�\��/�7�۪f�L�r�A+/>��~/��K����?1�tGƥ�L"2��>�9~k�l�Ը��Xc�≶=\�دγD�A����0�
N�
���Ula} ���$��ΌE���C���� ���r�B����Pg�i�WS �-;Se��]x�ǃ鄆�~P�bj:u[)i~�9�^�m�9aU_���܄�/9G!���%��|�l�YjE ����y�͊���q	���h�V�
D����ť�r�q��n�~�}!�JV��)2�F�4a�g��Q�NaNw~�W�(���6`:M�p4� Ǝ�Jt���o��6?���>i�O)�:�o�~��[������������~W�F�J��O)J�-���5��.����@I7Q�:+���$J��Q�3!Ok��/!��5s����<��R)��=�$$�s������W��A�-��< ����'�}��aJrd8k�B�F�ѝ������}�������m$z����}���æ �$o����
]l�5m�>��ҕC���-��U��?��OE��w	Vʠ��2@EQe	��aG����F���82�e	�;3J�;������MFl�t��^k��_�w�I��T�Y������e�>������eK1%�(���j�d��#�<�����S�ڥ���B�y�%e[��%��Å��&�3�:�%�u�#�=܌����Wټ�z!9w8.ɭ:йl�p�#��Y�`�Kmn�����[`���Vƌ^����C�{��8���Ċ���8�;͗�E%V�י���gP�܀ߋ�ne�IG�)��9W��g�t ������mn��kE��u`7<J?(ډ5����ǣ���[��oc_����N��4;FT�|�nf�-��W���ʗb���a�,���R�[xQl3jsn*>M��I�U �%��o�cm�=��;H���9���{�S7�O�8am"#}�����Au��&�ȮefPdm�wQ�f+�0�����LW�Ҽx�g��i-���g�?�K$�E��Ɠ]"�������1󛣦1fԶ���$���r��yzͲ-�*�[����f$�%]w�Ј�H�ᕺ�P�&l���9��G�3��#Kn*b ܈�,I (�� U8����n���H[GY����@�i��S�B����kkd��@l���;=���#�����h�24��s�T��W�@��!՞Y��d�Y�ڟ�	T�J�������0d��2<I��	K�Z27	A�Fc��7.*�wOYkcz�i��+o[��>3�՜/���~ϕ)���kw�����k%@���x+-���M?��"J�o���]�+���1�V�}p�.���Pf3g����c���w��f4%w��D�k��_�+�b/Il���@Y��fs{��!�(�v����k¢"M�u�.����>?�}S���L#��mp\��,ytZ���9Ւ%a*�NI��f� ��ABX��,�y]���塌Y�C����E
I*X���"��9R�iq�����?*%�	7��-�K0�d�"��/[w�ژ'i�읉-���Q�N}/*;+`=&?��s{vڸg����2�'�2_�]�F��/�~��!!�#(�NW[����,��9��c@M��]��ƾy��qP[n�8������6�̝���z?�B=ST���3�!� �=��Z��R'�ύ+O'��u���Ĥj+C3���j� 6�H�k���=jH1ӆg��j�;d�*U�݊�P}>Z�@3����qZ-M�*P�A�Y�i'['�D5-�U����r!� tEL��=���S�7��5�|z��B#���`��� �ʭ�0=��V}�6�5�u�F� ���
�d��uQ_ᨼ�ů�T���:F�9�6�Q���maM풝� 1'�K����f�s�O�_Z�`��=����Q'�����^;�fǹ�x��F�W%�:�J^D��g����{=ޯL�bS  v�~o�(���F4_��S����3��F�0���a?HR�|�䚆�)/l�xr3��)���@��8�55���5.���^d�ш�$+�KB�b�Iύ�~oc��d�fs�\��3Āo~���ay!L匤 #.�#*�6��p�T5�*'�qP<|���C���k�|UX��#������-�w��=2+%0�����rUꊾ����8z:�{�������@wTӸ�i��O��#~��-B�ӚE�"bc-m��z*�R�-�ؗ��d-E�q�sM��LY	G�.B=�����ל�C�2��fα[�[)~~��O�ݰ���lE�e������t����3�F�l
s+U����H���i�2^0U?�^H��84[Z��u�;��d�۲�U�R�}���p��*����\�?���-���%�!�$o>ށM��DZpj�z'�Z���3�F{�9����X�M�]!��7+��,Q �!�E�"���V*Zg+~/ ��@�~ׅ�PfEn巏��C�6\H:w���� ��8��ᕪ�hY@=a2}����C�Q�ST4��#.0�E��.br{d�����׮����N	i�~k�X��D��F��<����׈�K���]V�}N�4`��E�ui��A�������u��2<�`����ax}z���}��(f�N�8H#{�= XPe���)NH��Е����3DfQLN�e�m)ŧt'�ܪ�<+�BgS��k�8sF�N�c���P��C��}ުZI��T);���i� �})m��}&B��7�@�vx�5����Pq�����e��|y�J����1~��g�����׾�sUAr�U}��Mp�s�:���v�9Ɠh(�f�B�0X��#S��?ˤ�(���yn�6QO��.�ԯz��=",5Q��s&����,���!��.��g��U}��廖X3�;���p%��'����I.\G!�,&�	��.}��i%��cZ�F*, f�#;����⩜�r��@[���?!�A���/���@��yq$5��sp�Z���;5�@����qV�)�7�zu���N�ul��?�gz��2��U���7����h'h�17&��[���D���pQ\���"���1�$jbJ`j�RBWs�.�(��ϴ��>뀇zK��i*�H�g�/����~S�������6�=Q�.�a8�����z�ɒ�;�g#�W�Y*�3C��J��ݽ�O�z��_fB��E#�g[��Ia���?���["55�x��9l<����"򈛇�Ԑ,��q�Á�$�~i0��X�u2��<��/�����O9>�o�S������춼�L��}~T�脇����|����N|~���� ��U\�b��>/X
H�[dD�[6���yr� ��*�|͋�E��h��jS�E����v��mv�9���?ݚ���Z�#T/���0i��0�0B��t4�� uw�=cR@e�~.����>�G"��'�k��I�(~�ma�hr`�!�(�H��斞���[BƇAB�e8��"��k���e��s�(p	0�L�ж:�����L�1	� �`��;���u= �N&"�Y�? �SoV[�Y�1JN
�U��g�����+��Ű9�@��L�#eq}���o�b�$R��xyd���y�p�A�U��K�����m�}%7�f�R����U.��ӳ�'��B@֓�hc]��z�Lh�CUS�|�&�kJܸ���:"�兆��:��=���J]����	�S�y6薾������<qA�^C�FO��ob8F3F�Y���e�����F�r�^�^�,��ƫ|F��#�xYQ�ķ�� �ܰ{a�z�Y>��r��s[NJ�=�����yBG��3��=���Ƽ��{��5��xЗcG��2¬@�B���Aez0OԢ�Orf2@ Z�P�i��E'�4a4ҫyTT�v���'K���eL��K=1v~6�=�������E�m��x��<�fL;�5��(	3��ao?ד{�{f���� ��?u 5lR^=8��"�}k���h�wG��Zi=���~szd�L�L�I�D��ʌ�����0���� q����������Sf�%�6p]�W�qS�|?�0"��z�IL��=�f�hC+�EhM_���.�9UZ=�5�Y5�%�eq,�k|�ش�؁4X�4E`h����&�혪�֒��&P+Q����x#h�w�O�-Q��ɼ�W6鿠�Rp��axY7��V����<�\���SY�����LZ�/�K8��7�[�o �`SN�rx8H��x!�'L�U�{x}t��5/S�M������,] ����x��z4��I�ƹ�oQb�vc�<6�8���'>�I���x�bk�X��-���Q�-�h��>$*�;����m������	Q�.]'(t���'�E*ci�a2���Hɍ�Lv�ɲ�`Ŧ����"��o�����ְ�i��N�dp����5�_YSƕ����X��³ 3˽�tx����o}��T�r�K����(�G���|#]��t����78��b��qz�Q������\���$��d�Bv���`��S�%�Pp��5�$�^Ґl�Q���tK�a���V7z��g@�x�%�C���^6�)��;��(��D��Q�젛��x�gr5q��oIp�R
�^�D��E�k4'~�O<K��^���vG���0B����qxTR&�4b�Uΰ=m��0��5��7]B�U�����T��N��[m�;�&���i^w�)p|��A�ͧ ��u&Y2�a��B��Qo!R	��
ʂ����0���R�!�)h��V�X�B&aS�$mYq6��&চ?�D5"�
q���������$��":�@�bS�.�il�M�Ȍ���q�ϝ���l�w7�r���o�u��]�i��JHk�v	Tc��Y��v��ӕ��#���1W���<�D���ȝ�D��P�P��a�'��<�yo[�.���O>9����3�=�S��}�OT��6�W,<� �ej�=�,ɦccsP4��Bj+��u�6��q
�{�ڄ�Q~�b䘇�����-�Z���"�;;��Ŗ"+�j���3I�})"�_X�e�>��fa�q����	ϞQ���ۜ�
wB�@�⩠�*�����p��9����A� �����߭�	^�ch�g�f`Nq��D"X%h�Xb�.8�����C e��a��cţ�/�/4�nƈ
,>�A��Z�ȴ��&
trG���7C^���	�_���\���B}�[����# M��\��>eЃ�m��46ꗠL���"3^:7��2�e�������p�t-˶ǻ~�H�p�J��j�oG��0�!f��%���o/;���;~rG��ЈOv�����ݲ�����CP�Y>��OQ�e�|z�'G�����ÁKn�D;�%m�jtG��n'�m�"*EU}'0��?;�8�lYq�bQ^"NsO�zt�M	��p�2�C���pN"PB�*��8X�{�]˟�M̴}�lLE:�`�H(�\5e���63�c�̽�V��lu���IV��-�9�V�G=���ELH.K�h6��n�.G(/��|%�=3��� �t�v�%�u% ��5щAD��������LȺ�C06��L���k�2���� g\\��N���\�z�_:�0O����Fv��e;��D˸�%��a��#���"~��"�1�i�j�-�R
8\Iw����0=K��6�,:t�����`��]���8.[�m\�6Ig�r���jD��������z:{.R
��
C��W�;E}j���0��c��a��6�b{��i�'��i�س�w��+cp�yp���d�����Ӊy��tDL"sKwK�ّ��De�uW�˻ܬas1,�Ps���C;ٸP�~>򮷁�Uq Վ�#�q����7?�qu�`�(
�g>��������`�j�q�[m[���N�0'��#�&M�-��n:s�N��-���/ŕJO<�4��0~B�Ӆ$� W��у �5KA�i
�
:� ђ%EК�+TV�n�kL%��t	#�]��C�xlU�C%"�ö�Hum���؂��ﰜf��$X�\�m�7
xb�p����w仢�yzP�nw�A�(Yh�.�t_�W��FfW��eN�5�� ��q��_��B�!>��l	��}pg9�F��Z��?��E��_aM?�>K|ƖiD8B2?==i�ղ%�O  �n�X#�D����7��u�q�OZ��&xa!5w���w�.��`E��_������j�����4���ۣ!�RN�R8S_db��5*KdyRi�f���+��b4f���&j珜���!�cl�u�us���E-mO�|P65'[B���p�.�����?���a�7R�������$�]�L���sk��������m&J#5����k��-����� (G2� �����b�d�7������)C����ծ"b.�yʬxz ƋHҺ;�/	/��|٥I�_�DH�C�*�EF�q�zn�;4�5�dYV�A
�\i�ǒ���Y}cK�0����m�Y��T�O�@n�E�7�krCb��v���ꅬ�c6��[@S�iPc�*'~��L��P�LJ��N�׍���0��fA'��Pn�~����?u�P������$�^�������r�t�l>������e����a��%*˾��Jb3>\M�>\_H��Q��\�1Y@��A�[,�U�_r��BNg,�.{;1�4��_u�nWu�nݘ�"�ZQ����e���0_P���s��\�G�4�UD�^���r�
c���i4�~D�lFQ����oo��ʨi%��Bϙn��̇�{g��d\��-�3�C�X3	��Fah�P��SL|�?R��x��;=g%�K]o�XgHVR�E�S���+.��t�9 �H��%"c���Z|O*�z���i3�W{w_9��Q8S������4U�&��d䆨޲�K�Q��3�	���-���jRN3���ż���*'6`*
N)zḌM�b���Mؙ!������?��O�c֮"������yO;�����zLp'jk��tO��ӾW ���YO�r J���9a�l}O^J��ir|wC���^�]S�
�w�s}�:���y}٬�4ޏ����1e��}�IUy�c�Y��J�d�t��wQ��Xt?X���r�\�0@��.색��$�e���N3�n!E{C���ߺ:	Z�l���2��ܧnҦ�Gh�h�C��o/��F�YF��祣j�MU]D�ʔ�g	��CW	WQq3�I�ZƉ�*���"ER(V������f-�d��)5p�5>�a�u.`�܅�Ʉ_F���i�Ɠ\��3p����း8e����#�~6�9
J��3iN��a�(i0mG��8�G�XGi,�o0�f*>Tk���!ˈ3�!]�5�lG(n�P�ڪ����1D8�^q��+B_X�m�3��dC�\R/s��S� Dwe�6�/'�/�}[3������v��0��Eպ�q�X��P��� KU��ғ(�Y�:���'��wtT�m���'��P��z��vl�D�u*w1�[�.�E%�B�o�%�RV/C��b���WX�NS���)�8��I�$K�~I^y���X�RޢN��݁�Ư%�>��њ��r�	0E�n7�#E�	�����S#u	��rX����v$7�_�vBב�n&k�2zB�ڎ��`j�-�Ifk>.|�����MV����ɞ�>���-��U�8~t>�[�٩�7x��$tե$]�ƶhk��^�D.��¹��,�w��3�2 WK�͹��W����l�_+�P��t�����~R�� ٌ����
ד_fO�r���CN�C���Ѡ{�M�	�?��[⠷"T��>	���8M��� J	�
���F2��[��NhO�e���o;��DA� �0��a�����O��H�H�A P:���f\�.���*��X�/u>[M$iR�o�q��:Â�ڜ9A�ק��\��;q0���+��#|41�>A�4��)���)�_t#�q��c�
K�Z'��#�`��)���э��*����_�V�OA������,�ٓuOV����(��u��8��jRZ���Y+�:Py�)t�\�i#y32�c�8
���~I�^}�y�?�3q�yI� �O�\�����8*�2�O���� ����nq����SP�BfQO.�B��/ D�i����)F	�7p���H�ŉ�@|��z�^��2[gR�oo/�����6�ˈ�N�"��\"
e�M^��!:����-~v���.�Y�_1׋50�5zD��0���� ���'/|�:�I�w��tǰk�yX*�xq�ˈ�2-���Uu���0W]z���������_�'��q@���\�\��>���}���1�����|�[nO�;�k �v�aM�ے4<�˰�����s��69�?���r�����BW���62��y�-j�&��}j��������Ӊ3O�%׹�;�p NA^o���8�_� YٵY��w��Fr#�Qw#;��L��^1UEJc��ؠrQ�,��	w��(��bŶb���ʺ�q�hXa#l���n�JWeT5l6pI�$��h�	\�9j��Z�&�9_nA�@�f�F���E��v)�=M"�t� �U�\,��W��vDD�;��âdŗwB��hR趛[��j��x��Z�b���?4���}��5t|�jv�Ɩ��`Oi�Kl����}p'ȟ�j��K��Ց�\j5�֣���N>�3�3��˂�O!Iԧm,|u,�1��8�~f��;�qK@g2��2��B���<fd$G���C)�Wœ��Rat�Sj
dB��BT�W��$L��&EG�mm\��۞����쏤>a���	�A�Gh�>�t��{Y ���xċ��C�O�;Z��G�p���D�YU����;48�'R��/� ��׺�;�	 d&��g�X~K��KǕ�3B��K��z��w�{��p�����
��C9 =4"��\���ʉH�C'vHG�kznk9��Y��w���hλq���������$�Q�� L�<�tk'�[ώ�g�J��Cpe�_�{z�YLa״9��i��!@L�/�%y��^���Da����&�F�����˺w&�������v�ȭ���e����]����aSdlU�j���������cp���{��їG�qQ���qJ�D��|��u
���씢%�;��s��T�ѻ(��5�.bp��*�����F�*��@:b.xQ�k;�tel�(ay�DG�i�X�}>G�ϱ��T-�ٿNH�K�3E7��|&'��	�I=��g)�,&���ق��@�d|+���s��Des�C=��3��^r0��s��^5D���c��Pe��p<�����b��a��m�YD�/�%���t��C�VQ��iS�v�=5�[���$
h�U���0<�U3�����Xp�RfI,�{Zg5�	�a�t��^f��U��]h>���'����	AyޫET������1^�������P7�]�B _,��c��ZjX� �+��l�������"����&�籚� �B ���w'xkMFZ�����ꙖJ4Ǿ�P+��)N�y/\���û�[�J;ޛn����Q]��]��}�Y����)^j����&��ݤ�`�զ;����7��4�mX�(���j���ɲ�u7M֟yL���[���B�P��;������C�R.b[��u@n��sjOZzjS<��4��ɭ7�.����3j���@�\���k����o>u�|�'?pK+9�"��A$��u�{'�~��y%��k޸H�X����c۰����	����Pm�_ɮS�Y��c���(��D	���H�A?�H��z(��n��{��ʺ�ϸ����4Wc
��t�Ģ漡u��K�|����wC���Pv�yѤh��0��պ��r!��)-�I3�2���8�ڭ��I��I2�y�di�҇���g�����**83�|"��9�:�u�
:lEU�鄶��2u���q!%5/B��O,���ɢW�K4�1K���o��2k�W}ՒV�+��y/����X����g�6"��jy�:���RMɇ��SN%��P�*'�j�K�߷��{�¬5���އ��#��S��(�x)WW
�B&�ڰ��&-�&�>f��2�7��FtW��]��.5�ro�S��)�����'��nz���qK�i4�
�;<�P�J���k��.�����ic5������D�#��薐K��Z?�iX)i�R�q��Y%f��hb�8�׏�z�_��n�ݘx�G�0%�w!�y���@O���a�s��`L	o������s��%�ߊE'U����������'"��H�&BQ�!EΤ�t6�|�S ǲ�)�vV^����	94^H�ەļ3[lͥ_*�msA�i��Κ��^W+�'��З]��)h��ލ{J�(u�Yo�B${c͢8Tk
��؂���7�dCӜ��y���4�B��7)���41]_��<u��������3{`+�x������6v�Gϲ�7d�Կ�j�q���H��#x؁�dM��*��Խf�+]����4Mܫ�`?�/�};��x�\�h7����F#�3�Z(���֍��B�ٛyH���m{L��g�P��(̗�G�%^�M��f��+�'od���j�AxT4)2�e:4]�{��s���)v]7�ބ
=�	�7���Kx�3��٢Ǡ	,m� �$����&9K�>�ð�3sX�gI(~���C��.��"��tUt�0��3��l�]�x��5o�� +�+zm��,���԰�s2Cu�	i���9�|��D����C6\��	��e!�G��sr
j����и�M����V���xO,85t���sHc��k �+[�Yy�V.��~*��h�rr[��|�/��x��Kp�j)_��YO<�a��ښu��.[՞ߏ��'d���x:$Ĕ������WGl�٢�`���p�E���f�����҅�M���?7��H�q8z%��:]k���aʺ������5�k�].��';�^=���G��}3�B�.�9�f����)�����5��ͥ\�XVۭ+Y��|����[7�-2n,0�LK ��㤉g��Mb��V��~<^���Af,�3�	W1�VťSDH�&Qw��X�4�����W`�^/�+y��>��t����C5�Rʨ$�H���vbI�L���u,�+x�.�&�S�j�����	�p
,��U5�3+W1`]��P�pH=���Lg
jV>�0b�5����P��N��*���Mڒ~S�Uu>ܸS���鏐��
�1%����xxEM��[	���F6eȩ�}����@�M#��}��n�*H�	������0qN�@���t���
�o��̟��ޯ�w�����C���Kt�S�������<��r����}�3�d��)�s��Vx8�%7�2b-��pF
�븞r*�aw��߯t=�z�d�!�ww.��e��	�z2O���&!xTJ!��s�=�/T�p�.@�f�9���aO��a�lm�
�z�c2�t��F�S������� q����{F�ȕ]�N/�5kI4T�8f7D+j��o�*!�-�Y������Q�il=�G���C^�*6���h��rw'pR�v���R/5Ffֽ�B���c$�s�8����\>�,!�^.#g���.U�H:7uj��8`��y���,	�S�K8�����]�x�ڂA�8�4�ǂBYS��5y����������\;Y �I��X y�cu�e"K����tM���?}��TkrOٝ�1k�ʘ�\�&2h�v���9c��ˡ=����������^W��'���)�V�ܖ3��#/}s��<���~+쑮i�<UV��� 9k@���)\�d)*�ESի�������gtd/��C��H3�qN
ﺋ�&zk"\���P�բyd���*������8X�3Y~�V��S������]�<k�드ɩ�T���l�2��|��X���Y0�e+���t��k
�/���e������nP��pln!f�+�ץ��m�ŧ߅�a�j�֝_��6�$\�lfX^�}��y��c��l���-;i�ձy�2t��1x;����KBp
�����q^LԌ�*_��	gu��+�r8�:��=�V��l�u�dC7���c�2���i�\i�ZM�;^MX����^��_B�q�6�H�x ly���\���/Kګ�җ�3�D���ʔ����M�u��	��hσk�Ψ	k���n����_)�G�#��t�&!����Z"@����l�x��+��sAh�$�\i<���}N6Ϣ���-E��^,��܇�q���d�h�7X��Q㡎�
��>��Ӗ�!����W��ۨ/�u
�yŴ�^ߥ`�K�(��]&k����޼~��Ma�"�	$���{R'�����)9��C'j���ee��ql�=�Ɔ �#K|9���JG�ɃE��R�����dc�9{K�З��z���!����ŐtA��Ϝ�����Z��/����U��? Y����>��A����ł�?&�W���U�p_�"#h���M�G��!����ܒi�Ip�*�ʨ�,������-�����F�wI�j�S,R��f+���)��;x�nGl (	R�>�u.@�OY���d���q��Z����N���Xb�����JAڴ���4���S���ζ�Ѕ�C�Qb���KNm�zo��<�K�}~s7�
�*�ͤԮ&|T�g�2�������:�x�n����+���꟥"�Xx����
fL�d+�ə��./!7�Y���SX>��k��H$]U $�?����O'L:q��1�@E�2?`��ؼܩt��e�=�Ӕ,����t�w��j͘W|3��
ے��Ӣf�vA����`�6J��OWM��`J��@�j�/i8\�<h�"�Ӡ�@���G��S��g�3'
�.+�-#�q����Q�>��U
3�I�Q�"d����[�q8v`�O(���3��2|�b�.�q)�GSȵ�S��d���k�w�?�����5�������S�D�1��fzU�%�1����5��_��-�8�_�˚��!��%MT�g��.��O��)dt�y�t7�{S7i�wM�@�W�	��:/R"V^Y
~ir��P��$9"��o�(����7x����☌S��UI_�߻�Ɛ&;n�CK�ؤ�>�\��d���Q	bM��x���Z8� cP�4M����R��B�����0%�Oa�F����^y2ڱ�lN�>�kE��:ym׹�����3�U�D@&�c�s��%L���%�;�M�'ҰOCS����a�0��U�y�J[���B�Ɂ�<�#�.�j����/���h�-��l����m�u��|�X����s�vg5d/3�-�J`�"�ޠg�,M8F+Z���矧��o:�H�ѬC�����U=~;y�u�����9���e����Jy�w����s�p1愚k;�7�9:@-O?&V#���5r8i��ذ5x�+��#;�����{�C�_��vP,����[�L���+ƻt���1�u����X�l�yu�?�,ևs1/�q�j}xE��"���L�n��	_����I�a|聿/!�4����-&`IT�1��*}��.�/
>��E��&�Ur��~AL �_�(��@e�������,��Y)�{̢�O�,���L�ı�j�>�0���K��$�-�.j�-w��0o�����d���Li�@-�#byr�Y�e��_
a�@7���ZI��L'_�-�7�z���K�cd�cb/\w�p��A�mw\�N��n?����; �����ɟ|�j3�)(�q���uEY�Rm������=1�o`�y�p{�nU�s]� [���Y�G�a֮c��-2���J5��Q��g!��I�G!��!�B����5�**�yܓ�[��3��~P�Y�~�-`�r�.�`�3���֍C�{z�7ME�!56�������i^�	h�����T��ҴYs�aZ�\� �������C@2%����%)�"Q�^)��o�rI�;h� �>E���w�;��e�K��'��q�X����oO!�ض�S'����G���$C�Jd�g��,"�H�%�~�BxsV�h���c��4`��2O�wZ5h]bÈ�g^4��[��N�X��D�O�\{�k�޻u1]bb���KaWt#�5oڟ�y������?��2�����i��:���g�?ka������/ �
�09�W���#ϸk��M_Tf�I�f�;�-׉Π?/�m"�,W��kz��nwZ�[��	��<��l�.<�I�`>|��4e�ĘF��ѠL��u���ʭ����;|���򨞒f~q��>�����y2�'�r�?����tA+QΦ)�����{��(\���z�D.�̅<��մ��g�-���s�IE�Z]��y�l�v�	�C�_�6����8u��
!�Y`�CǇ�)S�5����H�B*^�Sȑ�d������vH�_g%!� �߇�����|{O�Gz�:s�|�Gf�/��j��ɪ�&b{I��2�̻Ȗ�F�bؽ����49B����7��~?a��ކnW��>x�xsEK7^��[�]�s,�,���TZ�3W�V��j�	 �
g�;ܚ{�)U���6"K���RJA�iد���Wl(��v]T�DX�h�q-y�q���_;'IM/�V� �}rǂ��0��|惫O"w���ao<$��1m M�5�8bt����I�=5^�q~��v��|�ЋKeq��?�4�D2����Y5���2%z��{�!�0�H]_��5��J���U��ǃ�\�,�� ��(?^�9��P��w< �4hYS�����5�)�kt�K�D��L����yg�=��ь�B�F��CaED�y �`�]k#ma�M�U��E���k��1'���6�K��M��
�f�a�ܒ�fw�72�b�S'r}g�8�m��֓=/��#/�їM����!]�Җ�@��5C
RH����QBJ�T<�U�{7��Z�b�L˓m����T�3��F�RP�q���*(ʽ��O졵��Vw}Ґ��XHB�I+�X?s��ř�l��0�D'.��6��)\������)�V9�U�s���~�=aK�q�:�Ն�[� �� �a/�D{j�,>�ѬRP�l��F�h#��,�~]vk|�4b�����30@�%� H)F��$r�$I#6�E�q:%�J?n�������	�i�=�N�� ��A��acc��Fj�����h�7)���*��J1;��Nc�*����3Gv;E�)���@��Ϩ+7���b�pn!�uG�*�h�9<�8`r��/����
��v��6m	(�6�������"�o���d��ζ�'�9�$L^^xp)�=���/ء%_���8�����mQ�vg��Q؛����C�L�:R��T�>�X͗�C��6���A�����S6�ܬɸ��;9Q��հ��Ĥ|�F�h��$p�jfS,��wR��V�D�h	�A|���CGb��iG}c�<G&��[&/�;��#� ���~��ܠ���w��6XJw+x8��˚�N��H�aڑ�b�)�! q�O��"�bNo�gm�$��O�#S�q�n�M�"���O���@>�Q��qK���������X���W��.��H;7[=9hi�\�f�>&T�S��d�Rv0�ұt�3���:����Q�-�wZ<E������^d����ؙ�<� ��nӛ�B��VwHD#9��<p𑃫�gv�@t�	�܎ތ*�*��[fu�AV]w��| �g�>�܌lݝ$��?bH���7��
XY��ޤ�r�`V�.��1@��l�������b�Fas���YWI���݂�!w���n���Վ�
�m������������-']2��z0�H��Lr�����B�ᗴ��ݡLn]�\i�9x��� ��3�u���5 ��
]J�O��҈U"d�C2��|
���-�mI�^�@R�hʹ��Jo�=�X�'W�,�����jH��ٔ�*	dC�P���t���2�~���]��q��O�M���V���'1H���Ϊ�^�5h�����'��F=1�η`�t0���b��ԕ�f�]��D>�D����cjl��9gаO"ψ"�OQn�ĺ[ጶ]ǭ�q!������2�XmA'�ԃz�,4�" l�b\�^7?�ξdL�E��U�(�q^�)1h� �L[��şڄ��`�'1n����'�W�y�e�RLv���r*���L��h���oU�����J'�?��hN֍
��R�A���Pl���=�XGX>��J��i]
�s�H��� [\��(&fߜ;��|D!]�hyw2a7>��e�9�/�]k#���M����$�b�����|����9K�S�õu���t�y�+AR�'�se��nE �9�) 2i�S�����y���5�[rK�	=�,�P�;�p�󀄵��	�>F��� ���f���0/��(ޯ	4����MqP��Sw��W DѺ�޺��Ut���}��(6�ȱ���WR.�W_hW�]n���뭾�DM�qȄ�*� o�n��~���O?�ē0��BKl;��(kzm^򣜍y�+�M������+'R�������c�G6��T#�*��:�z���s�P�{���B7����]�S�X�I�aPz�ڼ&`���i.��N�����DA3hgU�O�i�t$���]�ϠDp�o�o�1.у��?�[�O'�<	s�)�e����>��a6��h��V���WF��h#2;͂-p�㧴vFf���~�� �E�:�(��g�Ԡ� I?���!*�#���;X5�}�~������Q��`��lC:_���_�Q��
�x����A����6X3�������!�3�	�Y�J�v'��S��Ũ��¼������PT2|g��s�����-�2�.���'n�'�*�.GR�o��l9�+�&p�G	���k��`���c��*E)çOT��	�����v\]��r(���?��H�5���x�+�/sl�"d�	�i�
zκZ.	�F��x�ZD�r�?�=\T���/5]:��K�r"Żc��1�"L+����gGUCɿ��ݽ4���N�v��a'�}(�S��a���P������������ ��=�JA	�ޔZ��ܡ���8�l����W�2W�&�S�{�(�v=�p�����9'm�pŦFd���Tqz/�� ]c��V9����T�J��-���f�����O%�U�\���_���F}�����)X�2_�G�W �ڒF���D�Q��{�i�<\���M$�"zF�5�C6�Y�3>{�q|�-���ϛT���}��8�M/�I>/+�ô��cb�2���W�$�Ң���ܓ�K� 朦����(�;���q�1}?�)Xz��~�.4b=		�c�U��K�5�I\��7m���L%3,l�&IXZ�:!(�
.��BVdc�!���w+�!q�X0�� ���KG�8i�I�l�����_ɜ�U�|Z�|���(��ۣ.�O"\��������LS���W6�Z k����G�d��B����y��/��w
	�9S#��Buv��5-A���Ґ�Y�h���k�r(k��>�o>M�����H�v��|��d��otQ��`��L����]�{�g�R6gSY�z�Y��Y��enVi$Dde��M�S!,���¿"��vO�֫����|���:��_���2����0���G%_X�S1�q�r� �sB�lT�N��7w�4i'*&	!�j|�cɔ��W��p�����c��;�Ea���jlNf,#��@Y��Re�(^t>��U�ɦp�p����nE̓,1����,a9j�ۇ�ɳ�FO��a�紼�M���\�K8	A��cs�ꁒ}"_���f|������+	�35����1f�D"��S�\�Q>s��4�Ru���!�)�d��~�����.RzO�253Q�2)�
C����yp�����!G�͎���ZzI�g��H${��q�E�ݿ$$�v}����e3�R�<]5��Ƶ�/>�7���-����I��8�/MUt���L��+P-�]Ǔ�sޢ�1L�i_@�mI��^��Ag�7 Y%Ց4ܴ�N <���P�u�Bb���X=�*R`�?xs�Z��kH���Bv���'/z��3���@ZI@&�y� l�Z�G0&��\?��Ӟ�d���Xec��=w7,%��Cz��D���>EU��I!��yDf��,����9;�m�*S�;�o����ȯR�6���Pߖ��o�K;����t��qrI�}x�{�ú�k	��{fa1�jX�6i�e�S�E���jE����^�7p�RF���N9)э�����	�#�x��7$��%è�4�̯�Ӝ+����#};+�"���4��]�fn�g�����8��9�|Cv_�ۈY^f���\��l�h��TH"V����Jj�G7��m�@�����a���F^I����Ėf�u-��W�T�@R�
��i���L���!z�ZL"�%���:Vy6��.����w����j�; �Ж�@�����䵽:���/����p���H����A\�a�T:kEd�շt��&��w��4�I�h����._��a��S�~~�K��J\mg����L�+V�{s|�����w��TFk{x�m���g:�Dc���ʹ8b&�j�ح�� �T���$Fɷ�������{�M�o�1-���gp�	����4�d��D����m8V���D���'��as`֪~�g��Ƶ{��f��I2��є�$����f0�Z��l淒A u����bJg�|,`?�{�ήP�+k'g��g]��#�&2L0�(�&A���L ��n���};?����uY1ޒ�:���XG��=b�nP�$��TB��3��w��3n37��)
2���>�h��GS��	s��� =-��Xv��V</���|쪽hf��H�����ၞ���(1�;�fxn���|�F?7�g�;&M�e�^�O��bn�f|V���M�X�"����F���Ti���?8���7|*b�T� 9O�9T�75֌]�FG���8����R՛Ot�Y2���1$K�e4�0 j����,х��jc�~N���A�ŞQU��7<��hޣƚՍRR�{C3Q|�{��5ÈHף�<�s�:�=�f�t���^�&��Aw���ۂ��d�Ɵţ�r	G0Y������|�#���]�U������r"�r~��D^ԥ�C#0\���+���"K�������DĠ�Ι5d,e��0�f���M��fK����H��Y�Ă��Ҳt��V�N�p��](\�w˷��ܲ/�}�R:��SjH�M����b�,���3�3����;����U����g]#�D`�_�(ӟ�wDY?#�s ��2|���!��#�lu�E6� <��*؏�MIt"<㧅�����*�ΑP���L��Y�|S5�Y�����	`G��KQ'ث�)5|F��Y樵�^�z�ѥ�92�t�6[�w�lZD�rO���!�[P�>0�)��us��PmK��!�|���b���O�"��D�38+����i��F'Ŏ�Sm͆ǐڴgY����)H2�]M�w�Ç��]z@����1L�G�X�7|��څ���в	<��u�֦[pn�
?R���6���˙.��r.x�� Di��нH�ޫGE���?�p	sR���A6�<h��"���X	�w"L��Q�?=E�<%8-^��sI��>�h��4ཊ���NH��6�L�>���Sk��Z\�Xiy��p���9�@�N3:꠾3��G�Ƣ��=�K�r$a�X�6|QA蚼ߘ f)�|@�V�����F��[c9�Qg;^f�w�'Z�h��d�DWF���I�fթRI�Rˣ�ʸ���]lɊ��������ѼO��ą=�	)Q���`��.���_y�N�>'�J�j�w��G�:��SA~����d�@\�g0<}��W��b�}j�N/��=G�� ^Tj{	��N�Z�c��D���	���br��~�`��B�n�b�zc��x�LI~�߼�m�C`�G\���@Wr<�ॿ`8z�hP;_X��		�� 藬��\�n��?�<��/�_O�6B��0���#�bz�T�-踫3�F�A�<��?��)n,���?�У�����}�e��Ōs_cD�0x��V��+0�J5+�ғ�4{T�#��_&4Xw����h�iŴy��bf�=4���a�j�5����a ��o��Q���k�2dh#��bl3�sm���½�-棡9�[�ơk�3���gL^��V����C|�b�Ԑ-k����c����+N�PlC�ؐ
��~Rs�g.�)R�>N��y`>.�o��;q�b�
���	`Z;��:lkHˋh�"�L6�+⒎f'_�˥�:!����Ù��p>`cuu��'*;a�ܓ���1"�1��ao,b(��:�<<6-�<��҇���������ܪ�D^|���68i�{Y�
>_*b�ym��R����}z���M�)Cr���b�|x$��I{�������ߨs��63�*ڹ�L�� �/�W%���ۇ�[e�Z��Јo�%z���3e�n3�߾���<�
�t�g
 m59�9+�X6�8*�"騃��ȏ3����{C��p�g����<�x���N��ss�ޱ?z�����Uow��MB8~�(�q ؉?!�'+п�	�Q�9����������K2;O%�H���*,��c����|0u:^%Q��9OI�~�<��m�K;���:J��)[5JΕ�
��:���H��J�iDz�U�V8Ơ��'�{�@cMD�f�b���<�;\p�].�xi}c����_��߁K���뎁�Q��	XN�㯤�ޯyy놝g�R>�y(8}~�ݤe�.�qm�5��դf,)%�^V��,��?�j�H�|.����8��P{L���΂�����"��0��o��)��M��(��y,Q��?z��G���],X�T����A�08��*3��C��plR�9lӱGcÐ�Ӵ�#O��CO0h�r4�OX��b�C�T�d&|@���m��/�4��@+�X�P��s�\��/�3L�Ƞ�rb�K����nU"�V6����	�HZ����ŷf�m���T������^4أ4.���ޘˆ��by�,{+�9�4���:�F'-&�쀴P�q��d�-.�N%�οs�﫫ww�3s�C幁J5���+o�z�2�b�1��:��fs��l�&��S�o��ލ�v�ɡ�O�W��Z ���~'��«��u9�-������Y*�g�D��A��l�2��MgG�hT����J�m*��z�BT��*�[��0��R��*?�'?P/ct�8� n�il�1�U1��H~�kH��@�{M�}�������ڴ�ff}��J�j"����D.'~/eV��u�>�&�Y�_��ޮ����d���CMp�	#h���Au%�w�`jmjq50��}<%�Y%��h~��:5�|Z��
�#����:[A+@τ��""o�ukɼ��D8�[>��R\A�'�>Z�7g�kz��ѹ�"���G�腎lƦ%9��Z��:|Տ�쵾��e�u?�7I���J����@���àO���!O�p�Q�e�@���]~�lKg�~�ts�E����{Zج��	��XQU�w�zO��-f+'`��6V]��8�H���1�dO�t�r�,�O(/8 ѓ�I`�[���%�5*�d	�%��\ȟ�L_>LZuRZ ~2Y���O�L��׵b?%�����)s��2��
��щg���_����^���ωHy���ʴ�P�&�<"�����&;�늼����J46hV��]���;�]����
5ɪ2rt.���l)`p��d�2� hJa�b�d(L��)7������z�Xn��Y���-P퐪gt C"�f+��@�#H)Y�Z�(�pL�z�ڜ��K��Y�!�xŁq��u��2�p@��#�"�\i�J�4f�w�������g�0T+ûw����=E����\W�G8�'Z��!�f��D��Y��=}����Y�0]p�4N88JO��lҮ�<ƪ��_H���XD�p��ɖc�O�c�J��Q|�Ꙧ��JA@�Bm	.�hkzzZχ�
\Os^��,����C�05�І�j�:��n<`�:ˇ�`�Vb�"V��h&�_��<���ue=Ƕ���:���<rYڋK�l�J����9�Sۤt@T �v!z������}����Q��Ҥ�TV��?�b"⛠�`��P�&�1�Φ?r��ƛȅ�is��F��O����������:\@bW��bm�P,�lu\��|�e��-��H5DG5�)tG\�(}���+����8�����O�w��\�o�_Tdx �7�57C�JQ΃E�a))3��ȱY5�+aC�F�~�������,z����������l�)�w$�I�%
҆0A151�*���F�`7��}1�I֤{㬶�D���b�$�Yw�'�`;�K��C7�`���ͲK����k����T�%`0��Ł�m��:߹k��q��6VS������$�c`E�� ��M}vS��L�˾�i@���C=��v�{�9�6x\~[S6�A/�_��J���]a7|P�G�`H-�3P�=)�}v���#��ft�U��@z��d���0g�,u�ڰ�p��ö�iF��.�Y<��O�)�
��dh8Z�$� �PEFGh��Y\^�K6�i>��<�Y�JO��@69�l�獦��Un����r��4�n��1e/�=
tl�浹i:�;4	"���,2����#ʰ�>�^�`M�J���k��UJQf�H��no��Z�ʺ�'?�I�)��>�����?(�|�m�2�JY�R�m�l�8��5�����Fԑ�<�v���l�Ee-L��1�yJ	��֥!y�[�)�2V=ȯ���B��ϝ�[���>k��
".t�ig�tEB�}�ĩPE�|��9xㆌV
�,�5+q�x�)x��6��L5=��g�a+f��ݝ��u#���M���?���3��O���j��aΟ�	��Ͽ����d��F@��ၐ��]`�^�����QM��|K'��A>�w#�[�'��������ڞ�T'Y�x���U��'�^%[U�J~��nmz�Xn�F��W_�r��!�Z:$�)g��<�@N��ad�O��xx��Yk�V�'�.WZg}�u�� M�y�IN��M^/H*?�	��F�s��W#���7f%��c;�n�|x�t^r��]q#��h���R,����c�����f�M}$F8�w�J��:��
VQS��"IU���� S�5%��~�φŷ�M{�F5s�6����3hk�'�SZ����]N����#&n59�hB��5�U���v��O��*G� �K���6Z��@�^s�l�L�T\}�ɱ��<5ởr�ee���9�)�a	�p�FiQn�ƙ�y��8��\6iJ�ӎRM�4⩄[	�(0�U۩�)'ů�K;��X3�ݑ�T�}���p���?�[�1%JoC�Yt�s0kY��H�{�ԗ?q�K[����|�P0.F�+�p�����~���lD�����
��~�sp3��r����7����> PQ�!V�oUY@���]�M�q�y����͝�Hy�,'��e
цأW�:�]��0��/�Q��\B"���x(VH��a�8�S�8�}�ch��K5:�!O�ݩ��Y������bA ���׼ �2ÆYV?둓3�Sɪ�6�/V-�u��� ��Z.�j�؄������e^��Z��-��r�6L�a^r�j2�$9�cm��Z|b3l\�}s�Y��~?�_��������_�6p-����F�}i���h��v��uy\<�?��82���!>O��e��;�b�'��;U�!~	kBCc"�R&��#'���U�z8�?Gd W�����[(nD���da�̇�2^%���O��ɖ_ӁK?���j;�!�C��PL���u��B4�^��̑	�	s�)��r+�a�-z¬�(��7�@����e��]��3Z�ʝL�~��n�~�W9��`;������[�{]��^�%�8����l�U"�z"�S9��dWr����c �) v}��9�����B�=l�I���ٻჇB��g'�_`�4�8�ԩ��7��H��` �FZ� �����G"܀�.��I�~��x�̿�����ٲ��.���sU���e�W\Ό8k�ԓY�y��M������P���w��|B�Z:��d%�nÅK�=E����J��}t�!,k�����`,#��5ґ��3���*i^á�/�`�b]B�4��xV�����P=�h��2	G�^��C������������ɗ�[�o����ua������ft��=�$�%W�Rگ�ˎ�߈�M^5\���Faz	kzB�"�n���ȣ�-��������Xz��PtI^zPYH�,�ț$�L�HA��<=� `��.�,�����,k�Yַ9�dR�jm�б��w��:�A7���
���S�	C�`����YȧU�2܋0�RPy:��QYr�!�Q�s��MM!)��}=�f��[$�IF�I��m��̂���V~ ]�#(��H'�D= n�����W�i���`�t)�r��<��Φ��xܹ2���j�$�ZB���<*�t���V��=�-�֞7�.9R��pwX@��l����[R���n��΅��}o
d�F��p#v)�]��3������R�#%�9�Ԍߋ�1� ���{+�UF}d,y䑉�a��=��R��Si�t����#���<�4)�*1�-�~���KD(fa%�m��3��;Hy]#����JU�-j�b�jܝ%��i� ��2�t�[�3�Y�;)��A<7xf�h���j$�z{�فH4��h��_�����O����kj�?%M�.���u�k&���B����_��TA7cH��<��YL	�qi��C�?�`�.1�Ai+L),C�w_:�gR���� �������"D.�0�+��+��I�u]�6��d���e=�衣���h,���H����X�\.6�aGď��O�^- �+�#_�J��6.��a8g��CR��>8pd�~�~��
:��c�H����G0o�վ��UFl�-�2��34����R�S�����Q�x�� lJ�L2��7����#ئ��!Uِ��*������k�Q�:�m�{�G	�� S-D�0k[c��/:V?�,�����+�^��d�wb���zB�A���TO���0���̃-�My�3ֈk�C�����j��V)����_'Fȯ����7.'c�h��>?z�`YHX=����<K�*u���s�Ֆ�o�-J�Q��0�/�FF�g�s�?®�������m~"w�hg^*��(P���z�?d��P����{�x�B7�d�p�WO0�ѻ���}���ߖ�쵰Џ(;���l��@7���D-nhI���nk�og+��ϨUZ�q>���=�}�Q�@�v�=�Ȧ�e0¿�`c�[����e��+do���OA�_=J�cώ������q"�qDl(:��XF����S-�DۀU%��J�Ѿ��m��eؓ����-�MNLU�H\��p����]�(	��V�/���cXp]�uu���O�lf9�����5-t|I\���}��"lh�/�A�3\�>xB�Z������-NW�W��ia,70�
�j���UE�]/g�	��ż�'�S.�YC��츙80ϻ.7��}ݽ����n5�*��s�Mb#��G���0G�#��83�#�@���x���2�ZB�5����WgY���h%B��_���2FC[�LY�#yy�m���