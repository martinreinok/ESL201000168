// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
WxGId/rK4TNN5XME5rEkE1TI8zpJ8kkTlkCB24DDApQddTvXRqmSHCM0YeEKZ/mB
gSMMLXSIyHhHz/t0jn51xNN+0cMebM3nCGclo/j2ASKhUbVZmZEhd2/+5C7G7B6w
tOdsvwD1+Ob7FJR7UTr7AAoDX3iwciE/2W0KiTlflCAYPvv04Y7wTg==
//pragma protect end_key_block
//pragma protect digest_block
jvSLA6BbBlp76a50IhNgjiDatbM=
//pragma protect end_digest_block
//pragma protect data_block
XmuX7tB5rWHjhTHK7jsqPgPcnIN61NguTYy44iPGDS3M4VGRPpYJOGsmVA7Fv1mc
rGfjSgHKrj4l1n9cf2z+Sl/24x69SPuryfyHN/snkZCQ2MLWiHNeYufvaCDebncr
nw3fAs87QnqxNGSe9eFROg9utW2S2vEUBQV2IypVtYSqL/N+9AkZEp5V29gasg1J
TyB3n72Bt27I+66mnD7IobriNdZ9P0BVWnx/5RxC9hpdNG95gH+jOUrn1OM9wVa4
eu4czHN4o1fOX0jmH+paho6dCYfRcTBOu7pulBYBH89RItuxWNaRIuT19E4mXIgV
AyN3F3OGOYctS280cAM3+h3rfVumVd+yEWc3j2kzYLqi+OHyYtWxKri0IBuMIG5v
gQdDi58+/fbtrdQsqRdHvCrvuiyShNhwCXZCTsOeSRJHfaZc8nlaoVo9HajZq2x3
iQjuOQ90BrW6ZO4mIZu1/hQRd/JkArUOJ7DmgPpAPbtuwMm7UQ/9zMADFHIXxO80
OKdhPGSXVcmAyJXUUa0O28FiPmaBWdd2k6cKcNMSZszHYFfeuuSnkpQ0cP6Pfe/j
QEgb6ifEFkAKEEx6gBV1G4HzG5dmTiFKfw//IrWyNEHDZzVoBSGsX/5bNm3nO1Fv
AUVIJmECrFw0bft7K8uH3TI8EwXdfAan3ILlH9x4SGLTubgrUc7EaYHnNZOpBI5B
9P+xJ/HKEoWNWkFZ2ik6PI29ct0z9DnQalqk26ANZ/jBqfVNz0sQyJWcAVZtXUNA
Iff+yKDssqCwEjvY9r9ofmVenooFS8ahdddcisp7VHWgvouFkpaPRadzby9cZWJw
Gkh2zv62CMg4ZKzODfBXwUVL3YRiiozxsHr0CrIFMNQ+SdBkYb89v8Dd5AikEZJV
DfGxEGZn3+r3tnwFTgl20zvyxIUa9Ptb1TLfUIUSg8Xbm2pNvckeBFtW2vfcr2l/
MDBSb/K76svWxJ2RO9J/+whSxHaISqKvi/QxLMRfEaLpLIo2WHMs0qiuILCHnYOt
F9e6oFOvyll57q/MvdchKCXn15UqqRKOdC1POmCHsailPgmCEywF9k6pM8ww/xs/
t0nfMAXYXRnGNVz3zfKxC9XSl3yLnwymxJUyGTLmyVQ0Kj/+JLrYLOxy0KDuH8uk
ekswLLERboW6qwMnMuJqTcyb4MuLVo1Qg6gPDl8A9tfz1Gv4luzto1GDFIGaFWVa
xJ/Zss21DCoxSBKotQbwRr5WraO4hh8FbFxviMJLnYijRg8vVTs3V6oKKbnmuglS
/YH+n/ntWPfjlAXsmnvhPghNSQF18FI45qhna+saD9ROi6pXthe8q4iZz65i9rr1
O3Zu7+voAVvpI8rtPHO/2CLjKr9dpvX36aVI4SwGI9wuyJLbH8IeEGklzerAQ9GH
0gNI1lYfVPZl/YjM/iTw5XQWuqIVHfSE0Pv9aBwu7NS0eW26xOFiVWg39hvu0AMH
edgROiGmnaLdJu8uRt8x8YEq7E/R1AiG7HafBSv31J7Qe8Pe5Bi1v9t9cfXiuKQ2
xDFIA6Oqrh+zQWmHKY4eJeu3SuNWMQk/5uUKlXQnvPqOYui9TOi/1BvEn1LaEUYU
4ibsy9qeEHE0owoO3K3It6J5GKqzfNouKELA/b9s+3tnHuLUMmLYa8evlN5OOnWe
qUaIasGQkJBK0TVgjKGOe7ojTIR5qe4LtdEjqFjdQoD4ealKkOlypJwMZUaaQd/6
cMlbUi7x5rLLPRNuwKlQ4dT7EcugNK8NMDI44OXpsd+3SHMKTTWDsV6D9cDbuYEO
qkV3c/c6JV+/zIPl70X3OodrdQ8IsazpVFuyifZxzREnbg4hH/PSIV5jETSCEA4N
qvyf4Sn+uGDvOHLDfguvHxnleVE0tCQxBKh5jO7DVoZ6LFVhEva0fXVK1nCtxA6q
h6tf2rjvswEVBbuAWie2Q0xTQyI0bCE2L/KZ6wdc1/Pd5XoAp+t1QP5BhB9/j05m
NgsmDRqJW+u0ffm1scCTg7EeakXJImvRRPhzIsLJQQDgNQ5jfn5BiVgieq+iHuEA
sksOdpV9VxYaV+AOZuAAmQ2M9LS+RBlg2V1HxCFXw3kyhX9L+smWz4/IN+y5agzi
2Vm7w9+8M4aMB3Qv3c+QYzyClgyawV1JioCen6Eh8J4BKQ5XZZKnzU9oJTylqpYg
dVR1aoRo+YHM68HPsnFNmeanJKp0LgxomB52zE8hGiM5r0YXZFHVLQSnmI+yKQIf
z8kHhtZu8l3pCSAFwzEwwtbv8sVu3v4N8GaepkQkEbtBdqfhRmgi5Or19VBjccyP
iygRFmcaiyjcCy6woT+inZWhxTrdk7SVsuMeEtaEPIT13bb2+P6NlYhmAp9UKy+c
S/HlKDyXHXc1Wn9OnqYbBk5PjP2nwkWc6WaV/64j9FyC616fVnZL8NloneOcJ69t
zw/WRWIBt04RyJTCZNKTbAXQohWYO4uTUSgUboxcg516oraHei6oyW4EbkJmwggK
jkIygke2u7Od2r0h4Q9mUAEPVVP84z6Wx2J0ZeDZhhBP7ZnkuHSoXSgaieu94HJB
hqJL9L+NhruKPUu3/jg69r7+kLWHV1jclG4YWKayy3jSsybk1AiURb53XxC5M33J
F2fqgTtv2JBViwYFOvC7IsE2kDcbyuTpHI0DpPWh261F4/eIv5lQpcS2lOBaw9vc
9yNx+RggyBsT7YSaFVLchiveOiS3bh+Q0OiIKZ8ezkGOM1OYawpQJAftLmKVTCA1
4PFF8yzxj8hISEXyBkqJVVPMTuW7YXvCuUQ6r/iD3Y7Fhp25ZsdarOydGibUA+AL
VdCx7mFnjoLBuXtSwLkbYv6bp/fp7nRRPWpo4Jp2EEtKu1ar+ZNCMfpze2Nrgp7E
fv6A5ttTLTObCXn/fzlpMp4vKiQoOZcOh3g3pVSMnEPjBl0gqI4Q4Ibi60yonRF1
KKzwhTZzm+e8L9lgTzPLhJrjEg3MMJBRXFSxJEOwRPAKG9je9SN8+Yr8eqDIDlRw
dUKs9vU09Ubk6j0eplzj8PzJHCr/X4X3YAsaIvcup08CQfQNpsXrSsrUDBNpLDT9
NMElMdFGGJIzwIDZ194J7/JriWFeGzFj8uaUTzjpjohmT6gb2TqmlNhMmSCn7UXI
PNOSDxkkCy8qF/Zvygev7wCgZ0MboAa3D5L5OBG6H2Uh0hxePI+kE8fmSUR3/yrT
w6pdRtB0Ht1FuBDPlw1zAAKsY6n9c+/q5c6US8nL8Bwh3kAMsDu2PPUKbnwLh9dj
Ska1DfvolbCv7Rmjfany/B4K6mqoJTFdb9RoGWWtovw8tkIgvi2pAktmVIYwEHzr
EMdJaw5AHLZHxxmR0CsiW77FenPo/VtkzWS6jWcK0Lz2wnr0EObvADxjl11mS5TM
fpdhocYK61Nd/WV3LBTgfsRRNHDLgk4KLZpcIa4hkui2JCBJdfFIoB+KEBu3tHV2
zlfTy+9lHymTvlU6z6bw6U0qpnOUAtoYbHJ8Ec4fkjnZXBXRFBYvTuLyxfNhf+VY
nRwbIC/6YsTl+ABA8rgl7y+aU4JmlBRaMzcJp0MuUljN9WFcNKAAnmCw+vI3e2Yr
CXcRtAPHWXcxx+rOor7s6emZzhmgKEYaBU+AQseOOl1uqdozlNcItckBjIRFoWoa
UGlRoId4gU8asdLGkfFuIY+3hLDgVP7XU8ff6umEL6FLz7WcjfOWLYf9M8LgjD63
99JuziQsh1tOglIc31wL3tNOmTvSzgWbhAIDdq2/YxUh4jcTh9iWPbjd8n9xPO4Z
SuU9miUutb0vWhPmn9qiXiVh4NKUxHiUZ1ga916G+H3hrue5Dyf0frvaZNXWVTte
5wxMgQiI1D/3+CDaQTsrsWROn7zZMoAimPi9Xbv2QU2usiAXr2TsXFbFtgWiCu6Q
gR2x1opYf95yULhb2RHrJ81UYX4vJVkvl3irc1nhnTgO6ThBPmevPzA03q4+JHp3
p75cx9ZQZOT2zylw18ntBARjgT4zCc0dK38iJRhTHoU34gRAsUTv56UFTC9+U4aK
d06H+rHsgHqgPKxsmq1K4eGleNFPT991xuVDCNFB4pH+3V8APy8ZQ3hjGQ/fBce5
PfijdkM949/cibBXenUH3TsjUJUbH84X1K1F7P50I2E+gj+taZC3hiPd11Dvbjd9
k+izO2+NMNGYz7y1rP4zzp8UHkMqMhhsAI+3Q7PvKAHv3tGxTzdOC2ijF0Z/iXJ3
ggij9JbiYdpvB1tU7sMBieaepcVGz6vwnXYzhhS3y1nimwWnYeHa7/7aTVLe4CzK
PueIJMG6LTFrcHgcac1+CL/MdTnwf4yw13ci2v96gxqLns71e6nigcYL4TI7/iOs
oJA+2TfNjpcDTXzzssI7nvcnGsLohxG3eTGWpgrgsR0aV/xZk9WcN7anp92EX+u6
RTOzRkpf2L2mGI8a58AMXUh1hw4ISbIA6DKfXsZ0aZgRRLynIMhT0SoHiaHNTIjf
jCpgOgsRBSVVz343TV26ihkbRe1fUZY0cObjdF6sjfDo79TL4QayQNcrisiZrS2C
oeWgsm7EmLJy/eKSjQoFWBhHt7bZCEcsTqLkPJWr/VNiOTDGR0pYH6sLmbruyIsy
3qFBP9UfLgC2m8VVKWb7y3le9xkzJeWF9V7LJhYH0DJdVAWDqkV3OZtTqlmOn4wi
N4Dh+lRkXKybomRs2l1jHNbGi5HoN/MDTSwOh5pqBdgKrUXtCDb2LC6LHqfzaQIC
vgKkUwbgWl5T1jwV7G+iKzwu3ghhNJaHJbmDHKZMfO2GKtr1j47e7gD3HyxJ8lWb
PM3GMyzI2hIzKWq92nsgOBMIzyFHP78R+mEqDappIcnWOlXlXOzAvq9xMYI2bbGj
A/Z+vXJA/Zje5sLoK7wVrxCTsfocz6uWEayHM6NO9CNaoQ3AwT+eoZct5XvHfA/o
wDG//Ac5fXxdm9egkROQ+cOv0Ef5ynxeNrAC8ArX658a3pEV2fpk/kR7zR4W2NP1
+aqd9CZ9X94lteRk4AxloZuRllpAWov33wPjdef6MKGvIiEO/srDigmitCzQTqlT
jueSuuvcBuj6N97n2c59a2t850BAofi6gq3zqCMNFlFxIZJLnqewekgVkv2l7JxU
tvymR9AKjEmaNqhtC80RwKoaYTEeHMzHXoRZqR3GWskoWXiIuWrogXogs9M/w5fV
Aj9mP62IomZo+nb70o+BNUtX7xapnsDaa4ZP3xnjwcvjZQOhEG930posKeITifVs
XOfAgVuZd9ef9UNclgJRoBvelhaRsg63ux3GAghmxpmpFP4cXNCa8hP0qaMhcQu4
obhPvY36SmYr8/DxRo8QeMLD+LMzrcJJmqMd0xudv7vLfT6Nf3IKo1DAJPuj3aNi
hjYuNnLuDeKez5x8tSDaGowAunGS2QLuqQSX+uS8Ib6mOHeUh7zUGH5ckCCtMK/8
tg7dnnkVj87ktHwKq+8Ok9vBTCbge9r5x3zRegpxGegFQlJAPD0whQZa7tZ14GSN
jHkFJ5ktgVmQiqL2OzWzgllAZcaIvcl2zCxb4SF9V5+FTCLVX8DhzOCBH5K5pe5b
NIYq/zaxHIeHJYS8qMElCzaT7uP+9w8s3ETQNOTK4ejEfMcJM2eQvLlUQJYRKed7
/Q92QeYUAkEDsU+OydcefVh3NN1LD/i3pVvrZaF5n2JyhrUneIQGmoN99UAp9aZS
ucFSb1ZJ7NQbwFawb250Yf+rSrlze0px0h988UlbDbz4RU4JSROBW4pCTKvfobId
6Toqt7k0V81OYzHyWUa18AWib9JhSyRpBXQVXF8fuFLi3djxJ5c1tht/tnKwrvaQ
o5ZL3LjpjoleYTwm+O26fu0jzd4gGK45hv1bbXdLivC5b0+2XKl5JUU33rtT9sYc
pjf8dEfo5S1R9tVwj+wf7sQrwNZlrArYZimjLugwP9otzHn++WkUE/2FBzj+lqY0
Z8+Khatn48422IW8yr7y88ASfFNgrlsyTe6dNuq2vM2SCCU3NU5spfObvg2YC0J3
M2sVFbTlPoq1gzLm41oJwaFbOuDerg87KuXRChVBa7MeB+HmNDwPJ/caUDgfv4P2
E5Wz75pRA1LNPhyAh2U38YCYCVhAneGPaSE3hlMjYwlI9cOtuZbT2vpDqVRXDDHz
p/J/DzFWzAOqxehtVAtE0NLpRVnF6BGRpCJ4Sv6RpnyYKP1VSFykC1MiNDDQ0rvZ
sAPxBodNm5XeZ/Jmiiyv/vqIDi1spTpWcNanhmKJlzvpzqArwz5qeirayWw40xq5
Wqnl4SsGhFBsyPl0q7/qviSvYcWaqjA29Bu9x3BXQKbmuwL9LeBvrplv36B8RCBR
BjJQyDOn+VfQLy1dwAK0nyEXeJxeKTHuClY5q2pds5QbY+wxtKNTYvPPXQ6paXqa
1//ZBmzqpoEBZV9ukLpkoP3sDrBGFMMqNDTMkJCiZShXGtjsO9zyYGUlELQXYBt6
DxvX75oCNl3dQJ2z5UZ8MtwTenCIvarCrbWEBsmwdfVsNhVIMR3Bc8ZjSo/UiJpS
jVoMP0aIJ4RlxQQJMh2i6gpqOGiziMnq7ZNDNqvToppiwSiYy2MqrruNaGSM0474
Epr1qTTCqdhQfhAdWxLhUP/XlDl7uS7Ht8YJrI1uwrrNKTYrwz8KNfaVmtscLGZu
+SGMrjbyvQjpSHbaPg2i/zVDcAA3Dwn9/3NqDdx3sz7GvJG7PIAUT/NJYDdkE4OE
eo36MQmU5muz/noYgWuNKsVATkO3GjVtGmEwtRk5zOHuaF0CKyzCXYCMrDw/1YDD
NjZArFVtJqMepYIga64fjb8NW9iC4zKc2L94Oie4iqqy3+niDWvi2dfUxqjF3ig+
1rhMMmm5rtjlQkco4P01tyuZCqJVVMq16EnRszNu/cNW/eK80OkTRnXIdbnZ0chQ
VZnK0RMK+DFdQTurGMHVFTwtxb/5Ql7AyHv0C2gSL+jsYicil70PxaUjyLKsdJ8k
ERaOawZB5OxQ3zs+b8T8v9m1QNp96bA3HNK1AmFqsBOJmYejV6pW9BDot5dTBHTq
iRGZR64uwiQ2qzxQNCh8Ewd3wvZVjNi/RxIPEz4aZGAcY7HJap7hgcGsol36K3NT
ppkw449oeEHyjaBCMtsEm+2RYut+SsuJNZun3xwAJaB+a6WeAHMY6f2Gyc/98KSt
TtYa8lN6rBjFm3n3UKY68Rt7a16/IAuwUk03wzyicJWm5ClOhhMOcMMr4WKNhhMu
AV2K01Uwzmz2dykaar3HQ7rB4zejdIQEManda7XmcAw7PJb+48zv5ZmqBhWnV5mT
ncTztNq8EyG2uLc/x01di4XJWYzOqyPkczTV2b/Be7P/K9RiFbjBKnqjSKMO/38z
m2e604qig9lBb05y/OF74eMOHw7Yc1TKcmRgHKS9oUTCivpuKh5cWO4jJmLAMdC7
EUgI0daT9AyT7BxTW01VNASOUNiA46NevaHNSrpwOV64BxMGd80fQ/2jv/J1Be7y
tis/XbaVlquU226FgMzbpEDd/s2AOAjaG4uACw8XY4Qun1O+yQ1khVARKXx3LpAG
1Q1DnX8t+QBDaM9Xvcd3UvBF54hM1M68zGGQOaGQexWYYN54g+E42SERthhX4TU4
gdYLfICy/A3BaLmLtQmqX59k78xPw+NpnIfqymvfJ2P2GSgjmo5NkLkDMduB0SCg
pQ0Uuwm8f/vZdCfa5FCfEaKXq6iH3JEqMSwQJawW5JdBmBShO92iK4bylIYkJFj7
fQHWUcZMX+puSlrMO3nSrS7uXbv1tpFhR9mbh9AHvj/NILa0XMrujsLStYyoa5Yn
rvZpi32AtyovyMyuCdg9TMt34owR7HTvHkSC6ukieNao8kGnBU9yqnPaJYb4FtPB
EwIbXHdrCsDAfGWQKpLnjea0E0mYf9CWDKIGOW/PnVWVhXCNvnFcgytijKk4ssGS
P1rAG7cbsFzE1x7EVzJ08fdXMQfhEtdhasPJFrBnc6J0SU5j+RQHCfE/FBEDLAx7
fml73zUs5LyOWPVk+EJ2EHOxGT0jlLcmKEviSyvGbNkBK+rflEAii+myX6dyg8/G
2gUjCrzchx0W9jc7L71jW4Y7yWGXHu2Vb8YMh9I1TtoqDbjMo1scbIpo05wZx9ld
EVEufquTRKBn1VdeEJg/2oV/GU2lobpwZsApkzjqZCCb0XrPwVt5taRRD95Nw4Uk
DVxi/YEjoi4hfHZwVO2oQskccmq4As35Au+TwPhFv96s3Vw/9Uom6uibUeiL1M/g
jVmlD0PY2nytgkJrvjGabGk4XmbfiuC4odPLwTpEk/23KZAw8xrOJPECFTW7nj0b
bG/ssZs4urBxld4CstNUzsbrtQa5bfDnX5jS+9hkw33MnZrJ+jnITG0Hig8KVbSp
kAduRSIAwS/B+OprgAYQlZYSkoKjROBH+97zjFYjvNafUJs7c/64+KVENFqryuHm
2yaGLnxQPyvYoeicoJO0sAyriqGBwXhdK8rzjJ5A1kHjB/+lszn1+i1X6xwpOPY+
gmnjdogu7v3VTSSNVZ67Y9u8H6Pxo+iMRYGjeR2CO1iPvCVFBVV7lm4RQHTpMytG
OzUqlxZZIWQpjUcZ5zCmJ2qcoEt0yGQU19ybFS1+j4rAyC9Zu0wi2eKKjSp/dBAV
T+0S3XRIEPsi4Fdge8jTr3eRT0us4m/qEq64CQznjfNE5RQuASFirhgOfSi3X7Fq
fuWCA89lnrcb17J2eJAe2qL1kxMuK7Gz0C9ukltjFehRSPzEfGDqOadhMTm1k/Iy
z9MQZh3DVpZZoJWufi6F2a0YnM8uqOEcN92gppksp3xqp1lsPGggVOrppS1jElox
gzAK+l6PDPH1mUwrXEQicR5mBRgUuxghgQQFTqvhB/6rwB+7Nzg2SMfds4ZwhGCm
1lzBozDS06TFmKW7pzb87mSFZXv4XZ6BRWYWODwXZSiga+zNWgA6P2sxfZnOpSL9
rWsH1ifu355v/JD9tzphH3wCPKtLirUVCpF8HPGJxQiX+GIkVGwSKPH+fa5JVynz
gkHCidutZj3SPPE5p6fs5F+jF8Z4dEBJ1WkXiYodpGx39+NRZj0mEPn1GWtNY3Lm
/VaMt0y/k/i0xZmWH3znLUKTtLDuJK+UAGsmpNk0XnbbWYSTpkZ2ZmfGyYeq/8qy
sPDrvHWTGlJxx1eefhxhRpuV7sjglrnehneeQPjVkgoPUKQJ9E55+M7RGRZ3UgGH
JT4IS1Mf6iDDOzeQVCKA/pDeH7yJ4wXIQdTZocPByyhVdlX57IIgU8tb2qIPbdsz
Is0411exwUvd3csIRi0oLXNOHuawwvwVG8Ebwuf7rcfxhPkHdNZJpS7bIS6AoN8H
aR8q5PSFKkojRYNCisg4hI9CIHzasU5u+Kf6qPcLCXNT9qgrH/sPA7GQpCIkMlJL
hcFRXabXmOG+UMOSflRuwPgTa9sW6ymWCi3v4SaAdnx6p3zId5jMKNrmp7Vz/Agp
5xFp8N9ZtC0hJyIwsVbk6WAl7j3G5fWGhZPU2GxTeqoyVyPcU+4w/cQ9agdC1lRD
8Xnq37+te9AqoiwxKcvDvvLdftDs/GFATe6vZ+9aSCgRC7BNWZz7+JLkRYd+QzXR
WICxFLiwxu3jUbwEpjCfX0gNPMu6H0zRIjy8+X/mjq82DVE1bNnovm+33Zx9Rm2w
0/WsbJb6X5qoRXtNkF2uK5wMVky3rqZkKfD/xy8Yzz7OS6kRvhBP70wYUCoSdTDP
nMTifSxbcN7W8JJbpMDXyU3PsX/jTfm8e6CYNZYKCsz/fx47B/tG5WrnYpWjJ8jD
xA1FJ6l15YtOoRtLSKxfooUdFS2PRu0DumQKmjoYSbKlZe9480P4QCXCXI44Ehvy
JxjfCm40VM5dygZaF6GBAtgtc7pvMalb0WQNNCXhOrXz9Zts8Sh+ERBK50yd0+qA
D8DPFPH8C3VBmDEz5HPI/du+8+8lO7qN9/Odsnbzj1zrx0gem1gjRI0xujz9sWw3
zpNAKwz9Vj6fMzmAvlDEX13xIrlE55GRQCftln7tUo+LMhAOBgxLcZVxLBU0x6wQ
6QtXMtLwtYTruN78hTzcC2gGJfPz6GuxIlLcKBueqZVkAg/RSDLeSMnaVfWz+Z+V
6NtQ9kU27eqeKCWRL7WadTBXYIttXmwL3/Il12ZD63a8plhMJ3s54+WniF7JZEl7
pgYN8qVxOQ8zizZSW2TtxQ3MwLk7FY8PBRpAb7RRhqoyUxb82N583LPKThaJE+LK
aP3Sy65QjtQmts44aim7Fjr6O2LHDpouwZSXl6K6ZNniQde7qPqaDH+B0y/qULB5
ltQw1InO3T+AnP3/lk4Op1O68AjOtTqH79Z3oEeF0/ErZeXyfU+BX6ap5aKvqU6Q
+kwD2M9ZhlrpaZn1sDsCMEtq/65ETbnKPDmr40MhGP6tSwrqAU3d61IO7FcNvng8
3bbXJpkQVepEQz5/aWNuWM7YufO3DLD8akBGdt4uTakLZLVH63NgrcUKq4PWN4I9
6C9AATuMlS+b8Aty6d7JNMyVHUi5F+nBYMRjUwfKSor0BSSaT0hy3IVvBwGQhZFg
Iz7PCuWp1WYq5oYN1hFnXMNAxungly3nbqOKWmuUUE3IpZrBVaWvQXNrjv25isY/
VQili1Edqm+zh3hZSouLeL65r0bOP9PYTFmEGM2tkVVTuRYdxRt3TugtQYZnPWO7
qcN5swWEDMKYAiY9UyyyImlXU2tJyHyZVbP0rHwSGC3h4IKLhBzfF/hg4+5FVGbp
qvmQKISeTQbz49L1WDXiVkhtNnEKYXrX5fwUHp8a8ZbpG3TXTcIo3ZtID6CZ3wYl
5/Y8nY0z8u/Y9N4G9cdX1ZbzU4xo5aZpUSq9xY1PX2I54ZiGMkeTh5k9Y8Is0FeI
xYfzcwNonGzdM+a0y1DJkCVnQ/AEFeRNhgrDtrPukyzpkWdhl4doCCg7CLSsuO/k
3c/FoiaboxKmFpdQi1ckfpEyxC0kfz9oTRFpyvBkBSVfLmciVEga8w441J/OEU7F
2PCbyWDCdWaADVlSgZxC9RmkHqTbhcfL63IbiIJfADNWD9D9eDT3xFYMjKRqp8pT
lp2igg85Rlg6Ld08eMJCXYi5+brGMI42GY6/aF3aQ4FdvSLuLQ+t3Rzn1pB42g3I
CmXFbfbKP28gd49Hq3st2gMAgfT1WwykSaCXCjrCSISn/9+oH2TgwEPmWV8EO8hr
i5BvHuNiKMPhXoFX8wBJS9rvYBx1frwrlEqmR8s6e90G5vqcMOEgKkVmjr2z/g6i
fjrhbvuiSC48QOiqaAYPWQni+P2lsgUhQWYZsZD0g8qwHiC0zx6LmO+1SsgulL1G
dZvVhGEPeEr7Ld0XzVuDBgfbqDYv7Tk5kClumnFnJFTx0u18emQd+IgWvitZsdZU
CaR7GKPuiyZOIdeRK1F+NPyHz/zfObzey09MphwkgzhrE4VF37I8Mr79nFQS5hDp
kuKTmFyLzKqrO6JYXmI7/DQYcBhmr5GD2Z3DGnbpPLnSJ7x8GdwuZBwdH9IsChj2
TZhG05RnHwCLDMFPPmmdzK3AIIeIcmHi7C8UpE1R8RrWp7Q8kKq0A18C3OFE/+P/
S5e7qmDj4viwBAGKHZElBuLZCGT+owOm14+AmuWc51JLaiMX0eEcGxHZi4C/+U+p
Gg+4kbT9ckXna8ZpGSRFHUWZKCi1zZEXwrOjBcm+eKl7KX2o0syOSBwdQ5k1bfUi
BW8crrqHh+1ebzojL36X7wbHsNr3C01SiCXDDdrUK7X/lp+Fb/x+POE5KSildGnJ
YEkU968n4/+X1omrRnKVjvEL7T8PMpWV/dhP6UstIotOFv9vPR9JH+D+89atAgv8
FKi9M7TVYs3gg2rdvg2T+9VmHXdSM5S4VgZ/Dzf8mhGCp6/yZl8uCAtu8TzwTGPr
CferD3K77HMdJMiaREO4FudEZCTdkEbQ4ynqEvn5SUb22UDFfr6XH3wPz3fXEzzH
ijLE2kc9B6yGSWmCbS85xjeg1cAQ0Dx87oi1xl3pGzVhnMqQ50P+t8xXMm6y/2LC
qBAAS7HMsRgUW8EyXrFvA4sk0oyB/KlVMoBNEiTJ9clyF3EcDFH4OWyZFQqTJAE5
xj+g/hFp4fj/LatrxQ+ofSi2Wl1yeX1kSGLI8lVU9l2TW+kIB32LYdVqqYmDuaTi
IpO40uPcvuLHl/et9XvCxIh2zeT5+gjYma8D00C5rWmD6riEA8ksvJxcp+j2G7IC
ViruOvEJ9CLYhMhBUAPGpglFVNJSBR/Smh5J0p9ipH3NKSkMNWus8Fab9bdlX87V
xo6OhZzlRoJodcQCHqxWYte3R17EK2ccJkZGrGkt2nm4pZvt3htLGqOVrcUMcl2Y
vwQXjkjcrvnlG3SdUXphq5NLl9PM8qPUe6OV+xE9s+IX13+lH9aAbWpabeIMyA+N
OyL4Cyh0h+zNEE8CyHkH8EGle1KbmTVPNYPg/o/SyzD3dLYLDWrEMPEwtFG7eAtK
M8GVFn3bCHopXwF8WBCYBTAWJKcRJ44Crsmb04iK46XipOb7zmRPYMgowhGOulnP
NY52Mg6/OmaajJIClR3z3fBinazBARB+1bkk7n7721RspjdAB1+Xz3rvLBb4rx61
E4+Eoxa8sBtPX0Movvr4y0rW6spT5u5NyLvyVoflbfeB85GtK6+KgvwN5UuCsDS9
ulg7SSjFOhqH4wY6qm+gdcLZAgsu7azfA0pWwmQyEX//Xhjs5SVUXIo8SFECZPqh
mBrEmMFJmoxTcEqGkra4VUwK0tbKuabh+xrZaoG4HahdQbfYkfq251HlaLbRx7jc
xiCSoBU5+nIk/jkx4gKt0YWsspR+s+UAgui7OaKLHB9KbXfVOrVNAjJfBfG6h22k
7T6GYL1BjIRWQSrcWzbqL3w3/DQ4w3ycUfdNUA9ceW0l/S9ak/c/Cz5+tG4McqrF
HRM9D+Q4sLL1c6B+6FiMs6FuVF4hmQ3Xilar9lne7U7kQLZo55FhOcfTX5GnG6dc
FvsyLJNQYEf48RIdcjmwHfY1OZ44O8waYH97ilB9WGz6WsdWyeaPhVSuhKw7Falk
gnfXGlYH/dhUH6H+l09uhXDr+UgAoDXEHA8RqJfawDecAaCvm0bFr1enhK4DpPkO
zVF7/un0aS2Wo3XaaIvlmHEtMoU6dHPCiBYvV2ySPAFBx36UT400/XErAfS0Zw6+
8jk/vTR7ea9TL2++1LymJPTU2o2mjXzpUH5p6NgqEZiP2CqD5AG41PP/ljrfVci7
1YeuUGIw0eWUIOz3h3MeKkmwpqtGg+7HmHtVUFk7rx9ss05omVAyeJp5Oomo3I8N
LwbunqmUKaWYbgZx5ohu2TleFrlx9rtR+9EHJwV7+v24vQVXAnlEwdc+/K5058C1
UfPqXXfKBzUY2ieiXbSfam26dqb4x3+PPYdujOcZbENFmTIEEHVfGaRTPd8LusWG
HOezZoaeWdtDCSwZtLBjUt/yJpcnjAxZ+FCU/X+TXz5F45fnyvctBIAWNGKdK1pP
Ngt08mNvUDwMUfQUhclddCcueQ15yLKbk/GtIt82WBlP2KEiKSDYuU0NRj14A0+8
g6L2fq9JkihUMSCWC/mKGQMVUkVOMMcYR5PsdDNEc9rTkQNd39JKIE+bvz7cv9IG
2xhx0aWz09qEhYdns8iNaQtNS3ebuwvAhU7OMH8nr2VBfGVwAwzNBTk6xGiO2DGn
cWcsC1hODN0vqPd7dDY6jvFdUw+4Q4DKB5uxqwz5Nh095wRYfU2yc0bUM/99Av3M
IxYht/pJ7lHbnZMVtQOWcPygFZVVqVPz3NyNHh+pf4jfxXP+pzl9l6u9tdakN9d+
ASVdglbK+mhFgxw+qpK61tRGY+6nVbN70qdBim0ptNHtaB9hMnCUVgIjFiem7hTA
bSRRFa8bijYs64vnLF0iUHrLDl4SfkMqr7aLPVh9Eyy6XsDA0UpukAt1PyUiNVHt
QbGRWMbdHRUFQWS+SC9CTAO4iY5wBGhKJi5Is/GqY1BK5HTkJQjp3/5gMzSLnYiq
6N5X96hnJocMSvjd/BkJLBU6x1I7TEdU1LWBZQ5nDDFxCH1/DtQ20qNJLgQmvh60
XIa+uZdW0DSVX6PkXKX3ZYQJvtcHLE0Je5pZloKNWFigojc9Pl5QB36OEd/wFIE0
qmTjMBI3jD4Vdz8wGSR3RE3WP5JFBimhN+i1htz1S+c2TzYYjmw1T8ZHjp5kP5/i
R6KX4eIwPWz9g5YJxkYmY8M9DBomusjPGOmzft5uu87Fh2RwaHJqh/mUkTbdHNnr
ncuHKlFdU4F6ajP6qwhWhniT6olptMMOYt3X2r5tOIb077Mvn86VlFdFoZrUwE8U
j5OjN0kRMPQi1I0g6uIWn8wiM9Xprm/PS1tlNBWGT3ZrSvM60tRpjjKlkOCOXM10
K4QPXZl62oZupzZSRsQujYksRqCS89yiRAI6YBK4XvWXqQAH82Z3N2imwHLETKnO
l2TANorpPJIGvS2lPkk0G/hKITOCCftyS+Ktk3Zx05msVFFZDi7MVPu+qPUjOQR0
t/iEIM0GXQIHpjib/Bs2l8YXDiYJdoZlz535SbT+lK8M/1z1VVwnHli4xMkV0Q9i
xfirQK0Au4JKP7UB8QKVyxz6/51cnOuHRhzrNdiZcIHlaxShNYyGnkOeLRudFXpD
LRPlWFZ1liRFnu3vJnHvJScomupn8z6wTuFARNsxscTNrftRP7GGh/46GnNe0Dek
Li4UjgscjUkuxSrPdBTh4UkgpbZ6NfbofMwkRYXTuKXjMAvK8ef/GtmKxoqXT4eg
uCApVqFc6nCUo07vfEJ/VHGhYAEF57/zqiOD9YODBmM4AS9mxZW3/2UJL7cxusO6
V+4ayqQNKFBXM2w4qaSJzCz9hOwODEbwHXHuoSUCi4ZHuMWVu7HEvFuNg5jLB24V
UcolQbNsr2fAu/9JX7GI0V7YGJe2wFNpGBLWrjBniuRe9klO4FH9ZiaStEmWRQxJ
7Zq2XwZdoOwuIH6CLGO7fQrNxDxf8L/Vd0ZZsvM3HUhC1RUEiGSsxXCtAGPiJEnA
9QYUw2SNoQTVtPYiG1glXLiZou/3ywUM9Hbg+9QQQjwgC9XLbgVrqn7nxdCWA9JB
lGV3cmMvFxDKP6uMVz7FkvpmaOQazwye8SLeWLDcmWGVjulj7NhJFjRrN7VeesFN
rjcM1O8MVXgsmPfIrULEE4J1QtaxHM0YEDLs4qlTGRT7NtHfSUDPv8/3xlD0P/06
JP88HZHS8W72TRGDGJm8wAsIoVQ6ISkaoDLJzChPaMeU0T9F+F1tKqOwCaytnyAi
UiXyw/FZlXUIkt0DGgyznBQPSmquZ8vYm1Lt7DaHE3nViQFPKHWxMrENZXXbemah
aMhpt7ZEhln++WeAOvWGpFuJrVDwU2pgtgxqX3xAtSexWWNlHaSP+enKY73vsFGq
cEX9OxwGFtWb+zm2UytDd7pEqDHp/Zd+G3yGz+zvgBJBHzdP3DKImTQAcA8UInu5
ld1BSyPOFTJMCjRtgNy6fWpBSVHWROtR5zpRdoWPhPfXKVV0rQLgAtao4YtBSEQv
EOPIJVpZoK/aO/Wst7dGmznUQAj32W2J6ZKd/ePzLOr2hcrIWGhv3DPzy2PvbalO
gCDqBuPIt9PoXUlBs+SxJDkeDDzuXJt6lA6j0JvZH4OyV0FYR2TWd+S2w8jTT9JK
FmN9cH4eHIVpL8nE2ErbVTAernJ7ArXX9IhXpAC3f+JkrpnlbvUwKv1pVsIydu9p
TNtkEZfBKppeqQlgU31kLmFvE9D9Wp2oQ++oNjjZXhORiWoJAzVPzNOiHMZXhnWP
bgDb1trqQ+ZsS1G/qD7vfKNzwwEyfO5dWdCnhC1XKWHH2DqhVDFwcprcbSHs34PR
SovmXqd7Au9qGuYPQZlytxJO7WB8e3CMaSUESk1+RW5vRYezpPMHapcNYT3GjJFv
LV/kHVm+7fy1boivqXhHzwR6oDdmZvSes8I+T1FSFFL4bE8S6WRpFIPnk0iRHpyh
HC1nMzp0XQTAOkyyacI0y7EzDlS4TMOh/W5v1H5ubG5hjeuTc13TZgBgiuohJs2F
3+mzmopHZUz0rCyayfYONuXCg5rUc1Ji2lElnw2ToodQuIhuA/2NCjlkbXwN0FDM
yJTP2Ufy3PMd8afZ4J8MYf5s2sqxOCa0dlwILNwMvPvw8ZzPS+GSoORIYmIxNSK0
IQjrRpp6amtMMuGhR7856Jjm7f1SaiBhzMms7bHblz7eboSRMcYhCX0hXIFUGiv9
w7QPOLP3qyjI4o8O3YJqqeAARniFuo0ju9D6gENc8rAt9R1M5vOx9pprM1fwQ8WH
q05dq7grACWn0LUcZ23taT2MAycW1J++7MBTgz8rfS/LnjrPXoV+A2aCi6s+WILf
KzYEio6SuvpFyTNyA9GqT6g4M5A3bU2fM4uQQewLYcXB1emRuIrt/ot6z+gZOr76
mChOopfHgnUF5aaOpAMVNFyIPaS/8jJmH770Fflh4mWZyaBTQa3njTBwIoIKnmpE
/6dLuj/R0xNhk42eL1EuckhEJEWVsNLrNTt2bIyQvgKLsMeJoU7P5T0uMZk0itEi
QJJiT2H5CUNqYy+i1CgNT3TtVa1/XuY8xiAIzdinuK96Nj0gd4Kx9Nrb90tz5Goa
t5XLKmmNDiJKTg/4Yud+hsUUOLNvCSvi3mTl6yHY4URvL7/1r68kAY68kcnsQiBr
26Rhn6GEeY+MOgKMOMNuLrPqXBd33/1Ln/NkPwINDDy0FEe9Zrk4npHtvXSX8pNf
skf0cQWLdBbhWfrm1Kzsv64SVznucPgsfcmTZU9k795lFxEvmFQjQ2Y58QejB89X
WmaOYVvAew7aGl4khDYSx1uPfW7fCODLZOIvd+PjL8iyZx/FBQBUX62LYGDbm6yO
a1Nh+bECv0Cg7Z849PNRz5wuLoS8tLRHERcTBm7xBE1RtQuUJzYogD/0LheXADhp
FNQwmkdR8KSkQBj32h6HWj/SNSjiL+oqbAn56Pa0+rDix1+opgIjNPCHgH3z7xkz
idgKTcMAh41MVPFmiOCyviFo06PTGMRgpS5SA67XqWA9ii68C2Cq0FM4Mj6/1OjD
U1JtTloY5yWytoMU7fcWGFrJ3zZbSdgze1imV/ehyoYyrRTh11ZnxbRRnJ3qxnBg
/HEytNtdm8wFSac5Bh1u4FhjoN7k/eomtZuv0UI6U0BEw56W+o7ymiL8bRmH/TzY
DNKXoOW95CKJ6Sw/Y63UKg9SfW3NmBF/+Gg1YRXkMNIcQjpMvTl4M4UlNnYFcUs6
w2VwR9ZbH+IV+Qre4CRD+QZEwb1tKAqLNVI6/cad7sfNfeLi5Ea2B/68loCj4F8X
NjSskEyui3fKV8OT/asGzUCdZbXAWd9lh7wdq9KeyOfIXdfmVcd+/QNUGePPIEu7
EHyvRwvkHOepixsiK/jP0AxUPOFVW4/uNyaVz4Q2hoiFiOZuGGvrUso0LhZBo74H
hQFIIkFI0PzRBYYfUmqZ9+HFNcguPJLj8cc1tsQHj0pc5lAl6GGHPSGyXvm7tS20
or7fKH1nOWiSM3197dVDgYLKd/ozsECjTJG0VrDPfwn1lE2p6GYJ0hMU1PF//oXC
+XFJFi1mir6rFA2VBPZZshAATv1LHzEFPZDkk04RKdqRTuZQEuVm+D7iSyK2aTDi
HZWR5qEHY4vMQ1g0dUIJR+P+gXbDKODqiiYI6iNzQc4Fqu8w2K+XPTzDtmfVGjIN
QqWUOCV8UgXTyBPNCjHa5KAkeWO4THsldWQU5rK1hGbJLN3eVlXwLiPl4wIObylE
eOLqnfOtKUMTK2cAStmVncCdUhfHoTxDfI4HsxeTeOxrwcZP+cyx6naX3W74b1IU
mz8b82vZfI2OiriW/5Baaq+zyKXGxvBUEHyXgPdLxNA0d2EwivJexx/ngAOGKr2L
OOLcgqBPn7Y4OlL8zbyPuBfprbYK4bX5iBTNQaO/frabkTH5JYuhKOx6Qk8fCias
/SGT78K+B6hHQV7fZmLonOMZz6a+CKXkuEQ5ftbOUqEy2q5I8Sd9zje0Q7sIRwYd
MHvoLumXQPaFpbk97FkN/VB6BQMF9nz5uZ5+KzbbwW6Bbt8S2TDEnbZr0oOvKLq5
7oR5xpG6IwB8NXmALtKGInAK1qp+6XP9kAuzun9PXZ+Li2n638TTSmzkOSY99ulS
RuD9DF8X2CFuvZm8SFeLwE71TUtqFtquI8OFi/WeiJom1eTIi+8/gVdpADWiSTJS
mSXk/JcHEFSNCRQhqYvSAXWP9r7DGwEQgmeEw2l/b1MNYPRVmljZSU8EK3i4rS/3
S7K1gKTnPMXlfFobDAc0FAoJkneqLZ447J5HUUItjhfz4ISxL9fR/4DwNmC2Dm4L
zr4F6Sj5eR8yqciFqPbgKSMxgXV3UlBhuCdT+0zLTmTTG9KZ9IPqvT5dK8DQrxZj
iaPDKUZCviHohYlhXJJ12DJqp+dr5vCQVTm9vJVZT/qwVUrmVU+bw+WnQiMbNkKD
sxPwcTD2UmnMMphBNgYS9IhA7lvjpfvBPm1y7eQRLv0JkAmueGyptIy9E34RkcOL
RJE/AYPqIMr+nmnpIYOLocP5DnPBIa+Ph58WGB2G4TOL0/yQMHUGwPc+VWRdWbU/
+4/TT8J4vlG5I5XRskyW1/bFu0eeUlOfu5gQctQo1URs+U+HGlswVeke8LwhR2zk
R2qeO3STT0zwi0Z/2vwxs3eFYCwKrz9MsqZ2QGFvQZmG3zNAFDjMqNOJbMCnF/YD
dEhT9HT74a9oJTBoCFtSwKLtp5YOWHYmVEVQPam7xxbcsHATf9JgutZ04mxwNWcb
l13asuroTRgBdwbFSzgDurQSrK6GYRRb9o6mokCnDg/30ZKmNVehwST3GHQsCoR4
pzpIdf5MAFn51/kh49q8TD2iMex1HdOGm6y2sVPNYIT9NZ4XO2gadoD/sSEHt7xW
L3I1TJJYask7/SLa7Qmjaz3eIvtqpNwOaLf7/5qxbFk7CsNQMiqYImFEgRxZH8s5
e7Lfj1/YOJHk6/CHgI+0mw3pkaFGkr9758Qhfc3b3I3Q8XTpJVNCuW40PhO82/zT
xwjE6CPV5NSzCjA8UrO9eMhV2H8KxsMKvtucTom7DcQl9jFwT6+rKoyJmnSxq175
sUyvZyO5iAt+VZtVB6iRvitB39Z+NkEXCywsrv4aRm2Q30XDYdPQzBSuDS/Q43Ww
LVc49X4lTgMdWPzv1+C6/JEf7Gd1QA96xAntv0s2wm54TsuSVAWIEPj7xH0IwjpL
RDL/YWa0ND51XZHnEcC7C1MpSoGIHAyK+xEsFjA7g7cd4l72bovAnKktQMe6/ex+
3KQuT/dBUdXBxqyOy4BWkAnceZIpCZ/F0kV7rVUNx3Wf5p0zNq8qZKFnzYBi4m/v
FFrh6VelQQpArtSGqBMF5tLyYi2UfNhzd6Lqz2hk2qP9tbC4EVSXxMYwNJ05xer6
pipW/CGKaseYLThYc4Su3CYHVB9Ygv8qLwbuO4kQBTw2bbwBRTPUxi+rrgHom8Wc
2nt+/7zvlhJJb+FiYNR6dng7U58tHDxbGh30TSPp/oB/4KBZl2Kpi9oDGeyLMrHy
RO1yhW4DAcch4PNvk4VEYBZ5dumxLj2E8ak268ft3syZ5Q2ugVUiL3gBd7OG4LWe
nHDe94b+sJVUGoCI19lxu4JE5FJCmIwCd4slLYvo1PSld246lacx6d17fr2c0xpy
8PlIeRTsV4EczIWmxTGPycF2A1LWJ+jRoSBlgLBoUPp31ONqSqADaDRPrhjecbXh
q4h+anlLl1qCpAMxl/s4xyOiqy06XhYrPj39UVKMzh/iKGGQ50+Lx95U+HpuKjEP
OGYufyQi8GjEoUol0WnUX7cvWUYXp5dg1dNWGgRwJIOzVot1xddEGBmhq4Aw09Vy
qVSDCm5KYV7tC7XMeJ+hhkZnjW/fX682LqaCdzPyR+QkzXNd7AA5vk5TMz9/U8tt
6H9jxmZF/Rk9gQHcZlsHVR+VhQD7eFuwznfD+nTSg6kzXpQQi5UQPMx4UoTiwbIj
ySPrO3zCEDWnDTerQKO+2BT4su/h/tYxynm2WXsI4xR/UdQ0jO0krLlojKwQzEtZ
IAPO30lA/kRj5huKzXebKYEv2g7vLX5J8GanKSRjiHZc7O5pTjcnTkf/rHb5ouza
03emhRX8W+gOZ0y4KYSEeyI2MY59lXghSdPZ+5jUxPC4EHQHwvXjwQWgaV3rkgwC
y9FRqntAbmJYrqAagEnxB2aPsGwNwDFOlH3sr+JYuSdWiuHprgeutlel0djI35Gs
nbWTiuqKKneYMnZFdleWB6em++i/F/lXNojdy3DbF4/0HwT8VrZ6qJqLq6RYwv+P
9i+mLxnRAX3sMrXGB6wCaU3TfqaKM3epK8WtXAXoJslguw71cncmqdsJ+GjL5EzX
RLFDrXJThoT4w4A9IMBXbRmGKJU9niKPTLJWl0bikGRjVpSVSGqzjhx2ImGtj9uB
pvIHpAJZy2Gtn+lHq7xTikg+hmp66rcZC1hCEcHw2qFf4eaP6sNc99mwXw20TjOw
vOn0gMQzusIfhAxG9UYHrsTNUUPbnLwBI3I6YvExCTPc6jura9rVNdyuPgJkcuHx
fz3C7DHQIPwMPtBs7ygV9nT/+qrr+zpZVQ/h1zs0d/qFEP0XUcAwV8jhPZOrN0YW
yDbh2bsjlyqgfaQBl4gxuIGuBbTMEUXh/tM0SdUPKTjYlBb+9ri9eEHaKlW9nLHG
DAUkk31pPoJKjbDNrilRKsO+3JHqYRLT+v5LX2d90aNiPxACxBd6jjxZCJRAHcJf
iddiuLYBnDer09dq4+lJiOauKRqW/9AB6As4ZSHo2TaJpriecNC9leygUXg+TBbE
ke1T/5eCI3fMw9MjGZTE9kzzfhFja/2lcI4/ENhQPbjERhIUoSpck9vejBmK/jEy
eIYnGQj4B7mAiIXIRUDDmzkeleRQseTn+CYgQkN83dxAzvBy+/JDnSM/v73nYQV2
PGa+4AtbPlWWj+vcu5ao7OcN6EhAba34tnUPshuAzLhkNhkloXxRvOwASuwSSPAq
fvK7JqRnPW8QgCxsTKct8Ka+Cduwh2bBdMKg+orFv1U4+IN7485YjegAUiOkiQdq
+71G87fBJmMASsU5Zv9+E03xirEayy4zfXBv6lTxyoEJ+7/mNxVZtbp7xUzPVkI6
/b3fhq63+zw+Itey8IyI1EDaP8u62ZXELxCW4QJ1xnQFnGjRkIxKWysSbIkOaD2w
7AOmDZRLkSEyt8ZdW65MQxiMCmvKoMMcXenwdv++/AxFXHr5tjWbZmQtJhiw0wTE
3VJtQfubIDXkZ8LCL7MiXlsxr0nmm0DbuW2mXcyDCLLvVEfSUr4EJiTGm7USQhs/
9AHS36SLhhWhAB5RPW3yzAgiv1/1gRdDwVXary+0OovN6eXv/IYS1G/Xa4uW/cqa
kHwxYbGlq964TJzK8Gql2z9vN2Kipci3z41aIkqZF/zCNxTGTKYgtIm0hz0tY3cp
y6IE4Xd4HElKlK9bnd658H2q6nPK6wg525+NDg9g8dYTV/t6iTXl1fo6kE+B71Od
IHyjcHNagpM1JJJkaqM5+RsJPjf1hdIlmLHaWPzuJbnh7CM+sVDWLE23I4VyXurX
jABDaKB84hhVhMI4nmBxQjrylbg67kseGPEKMJufSQxIS+YQkMOuFPiT+ABmlPvY
KsChf8fxnpNGNRZCY0XStHWBj7TneIxVKhnpyCnc+Zze0CsfMxG6qgG+u1yBaF35
AVyW7DWVmYAx05spRhsK3K1+yYZt2Jh6/PZ7MmSS0iy7KpLRhLxeeFDo9+Ag4zCp
MrSR99vyLzk6vCzNgRDWjExjy8p8ahKjp8fCqWXO/ieaLFjs0bts8i45a9TC5EHu
jgpdzPpa4ATVpdThfPCjTGprTB5B/MFpHsTJjFUfLL4pAtfyCJemGKZPwr+zFWPL
YsGNIqyJOBaSuDG1NBQOVhJfND6WtoPOf5aMcSAaPKyTsvOMAYmobeWdeRMLuJe5
HJClqEOEvG9pL8FD+DtMOW7w5JHibDcvlIQ5hTk9JdMc71TNBvznuhtnGVoBoUPO
9HitoPvZDpQymy8muz0lEuU+cj1RmYW6+ASy8eSGAZl+BA979ghtgPBNiUHTgg8J
te8MAcDInNNuhAJq/Lrb64wWrNj2/fgReTZ3IT15+pInPLcq8KWOYrNDapfOKPo7
uWINrCNYvYDlFJ5WqQS51vj63VRVggUyOomrvms7XCQdpSoDuc38oaS6dVl+rWJo
Mr0QAiVdVoQzliMgTY6wy3qpA7dG139GSkGMHBsGe79w4117/Bpk2d9PS6Cht2Rl
vv3qDxfgY7RhcCOjmq8lE54lkN1+EsEO2d+soJ/m7DnIG/+JCxry3cyX9Kr+t5sS
ScXKVLdIxI3AT+OW/fgZJwr3sCgDyrT5vNJef9pqMDj9HaPt992wTAN4tAcIQ6p+
vFlwZnLqWjx2AHxCYX7B5f2zViR3pyqbl0PQSNc5ppRT7UvX5gLkwoDyHKnXT4bZ
JbVgsLNzj09UdKw3Vn/MlWlIo98MyTvt7wUdu3ivhmFvQ8ubS87qZxMb/rQ41rtF
vyRB3kZHzEKBkt/VV7HwmvZPwjkivHn2B3HWIveo5gisEHt/UyutKGJDIIfxmXAV
mPhTVnkl/gzUJRP1KobIRj+nSMvVrEk7F6Ue5PYUxB2RalmcAufBliSSgsiaIdCU
/xXLOBIC+X6pMWxvHf8ko2cUCRq0oAviD2qJFwy4SPVVQ6F3K2zLUwH1Tfm7Q7cx
A3+xH0WQHK7HvguDf0fQUUdc/mknd+fPiUDlqoGaTHBWF6oGYoM1fhaXIMQugiJ6
MNtomX7U8VR44znkGfwOPFNCvMdcehLV9sjk87FZbeRf/dxDhHguVW3tYVdluTwv
02aWVGEKZUYe91pouSspop2pNSKO7E49EiZ6k5CXdRUE5h3V6OJom8MhVHCHfGhO
ck/55irIu+L1RtTTERl/nO7mqzvr7gItQq0AWy8FcaYKgp8gWdAWdELL0zR/R2eh
UZ8AfJOjoA03JkLcekBkHMXVraKeSn1KQU502E3YCEDrWudE4Rqu5RYYFEgFZsNp
IPEOhSKj+ywkjwzbDW7bADkQQ2keuwcO+EWGp3cthcbYs5F84OlKn952snEqhwPJ
6iVLxHjrt9Ea1S3snxMeHlkEl+vxwBvuHRoT5nbmE+LTUHtupJiAeR9+o7lsIyxf
lrpgUnwNNCojzgNUNRBeav/sG2P0pnonbIKwVO6OzGpDHHtOL9nujryivoU2ufJG
+5Xvw5EUm2RGACuuT/PaUJ5bVWVx5934lP3zERs4+lzKGQ/nbZoNcaP0Y9XTIB8s
JoOGEnYUjCvN8+z+kwe+gr6nOWyXuUT/h0oBN3I85La/skJ8m8YIy473/5vij1xG
8DRzeMTL42OliVLQnKcaT752MLL6V88wrICBrL75Kkql2Hh8ZlpJ0hCY/lMJF2DJ
IeWFlFo0kmfVaLr2cECbm7eBT259pjghpkiDhTUMJamcCwqmejo6mNFOxtj0al3d
7qPJsHTCvb6VvZRTcai2tM4w7JmhuS83r1O06rtvPrA5ShOVRwvEYPFXJHKQjcNU
JKRnw/hksDeSeQ/czBn72Z7d2Tmc9oO+uHo0vyBgL8RKldCGw9bZtVe464Ju2aWK
ULYhXvOh85c0v+JsN/T1KvN6mtAOV/XhcGW0hNn/HhWeYkRLqFXLyVKF3xjmHYVR
rUt1XkmLknFX/pu/eaxF2R5x/EJEIIcHDz7YI93rEV67aRVl1YH6WEcQRhvesLk9
OAPxj4xyWuetPcftEIy1P16fx7xBAN5SIzx3PyiTyMJjyommeMvpDfvJ8sXQu1Ty
dpesC3RoM3criBkX9EJP+FwYa8mxmBKBkzffr+SnOJT6o4G9TfW9sQYb5feo7kXm
Uv4iKHRG5yMsxe05OaglOlXu+WacjXED+eW8NSpoPK7H3lI8Wv8umy2A8S+o7Zlc
mtA1l9r4gGSe/BBFDALxgJwe3MChnzjESnr54279cIoDjKNIvW01DWhnrYp7g9s0
Y3ua9Fw0HZY2QGBqDsQTJJwMCgJEiHb2ivJiAKorqswE+63bUFW6lfE3fkC3tHQG
WYJUWzOoz5dFF7PdxiVIt1aYeuw0PT6JrB8sVEmFywL/GCtf3bDh1NEwmE1V/DJj
MFjVOlotF8tWt6HwPDsX6cfWKOE65bRl72/Q0uIbWshEVWtkKNmGzJ6p6Qz4ps26
KnAOdSdIoO4mOsl3IJu8+dO6d4F+oQn5OWSnMVvEyPVo+ftPyLMPrGPk2r/RGPcj
pZcXP9WoEQBdX8gWSxaPnygCM+RFcd+7h33FCIXLPk42lBQ5Hxn9i2X85DB7t572
jq+n0B+wrLz2FXeroNu9V2jxxSP7GdTPAmheW17NMi+X4GKgXSQ1rq3dmM03JQ1j
0k7FTNYailckLFRp1iZ9yMsDy7357zVLD/1rA6SHU/hHIl0ScT773gAtkzIiGDlV
h2U7Y9jpJwrKdi/RU+3i1uXpWiXlFdUu7FIDVTUPMUcSGJwtwXkdfHZzXyNBo20w
tblzFkk0ea20HofMwg4iTVlnwoFbaLlRbRKEfh/SLNXh+lfE6e/SEpYVOYYPUZy0
f4RP+blQBOcHpab/8+AqcoMavIbJXK6BsS00ofg/ycc0RgkTdjEmjVNo7ITcKW4X
xUF8bCw3AKEfbgBPUYb5iTtnc4q51EmU91DOeCOV01nOmYjENgQpTRbI/QlTyN17
cB6muAbzOXApXk3QXKp0Fy2GVE0XtN6b1s3AW7bX/yhxkSLYImU0nKDbGy5yLQuD
TiwPr+mU8xuAc4SvjTelwItnjyu3uc418caMzNj/hKIoe38k0iW2+iUniUjVB/8H
MOEG0GIkS8gaJOpmmY24nKGIBhjYriUFNYiBlym3GA12HyzxMk0fcD2QF/o0wcsf
5cfCzSWONImvwutDWcFM2xYS4sQeWZU6gMgnnOh8+EifkSGj0qRNLepRSBQ+2zbp
vbK2PNtAnZB1X6+97+gnIXh3KNfq26SFQ9LTF3Wg/9jHlEXF5rEqJQb7WHwAFKxl
u4RQapJolUjY+0Lz5N7gvhiY474qAFtOyORzCSPwWv90th0avs2RWQ/N9LccxQge
G2vgfbNfjg9XfladFzrdCDmggH7yAq3y416J2JVceUPOiYEEAdpLEDiEisNwGhct
7XmVN6LVcQleiKQp16rXKrJRR7ohhtbpMLqqdF8e9BI2hBIjbqqdhUOFb8qw0qd+
u+dBQYVlV52aRrHWkxxWogVJC0Km1g96p4PCJd2ceuXCPzLnovk5CSV2069GsTKU
XvHqurtc1mWo/F/zc6dFh4MLoII3NYXFWmO0MLDQhMW4Em0bban+e6NmCy34+arS
lPzkkE+UFsRXtvErkbUGwCpY+jUNzF1BBoXzfAlvhPb7osIPTXJiRo5H4BCfma3i
WNo7CZaejMkThl6bwwGPkQtwm9C9A9Z7LGw9jMTAFA000a0ieUqar7ZyZsHWsBRb
QVPoLNftSEc82NUU3Jx+pjvRBTDu+qkaupnV00Ne4xuw4cr1gKQCfAGYlYAl2U19
N2wlVEnrizarJvcMvSfJxYghShI+VBYkyblwtWTyH1wW+Cl5NgOderbAqHPEvk5w
5WobnHqqnhgAxMPcF6KgOeGvzccIGfs1yzYyv4pfy7ALc69gIYRlFTlbvMcEGgAJ
pXxB8gIYRaaJFGMWfuZNeB0bd3mT3X7WOuk9KoSfWmIdEJ7m8sWIZNmxFJH2bi8+
ig78CG4MJbkE/0uRow9czmvFAA3RToXFVbxss/p7AEbg5xQj9XiM8ANIxqVZVlbk
wIyMRYDjRd7eCqVxyODOQxW+iLTeUUpyCJGwEM5ZM3eiHg/xEabMxagp74e5EhEE
26IucVx1Vw5NlrFvDL6YuxmGoz59NdtNrZF6cicKpcssBprRQOfPopypEFlxM89N
x4AF2jjiRQBETBJQUifZq+f4gbvrNvArZwfMglF6rsGDN6gcry5GILznOJzSTKFU
Lk8KaQbS7GQUZxbIKY1Nni8WMhHUBeKQ0NmCrf6WkEYIygfpYEC1QKVDiNumBH/Q
h/ZPog3gCpke9p1yr04dL0XfkJQCXnmFamUyorF1C8/mHxzafNIP+plguXhMJ9vX
7HSkrN0+9ZweQ73xHMf3NC5qr5WMuerfve4JXHiQr5V+psUofVoTcXHrVSomR7uL
JAtAtg1nHPeZj8WEBbyCn00zuYU2+dJuULfKfRue/u7ZlasGc4EsZlYEgetnxEEB
9Hvg2/jgo5MCevxxWfLWHs6nISiSD12bOAgt70lY8vm8f3M6+rYyPJC40Phak8zj
wKXOkY2sChSvjN+fWnliahnJsxOfIwW+2EwyarDna5jMwuq34r8vpcCy3II5Hsye
YJNQiM+E0xAiKMpnHL+RIyvE9pSwrX4FILY9WVY0m171zVUL7j/XO5f4L+3eKCOt
Xtg+gOsvlfqNYgtQ+5y2UDN02OR7QQ39GFD9I0DNfXioLONktgq7bebrdgwD1txp
371sqd8AG+bihDUnxoS094j3noy14C4waQoIDM1Hv1Xiv4ky8glDjijIuElTAJ6p
f1BCUfqLwtoYO6aMxcHKDYFR+t+ipMGpun6i+kgZx+wo/Tp4Lj6FoH4+QjsEtv/8
tvhrwmx/kaBq3Gqfh4bH3TUcoPeBDhB6P4b68vd4XKeNeqr34uckiyDm3LafvKCl
3MUcc49znTawmQb2jqTVpQKy4XzlHS8STK7cWF6EnGSbjAAsOLVcN5B6+ZUd1SYN
gDtj7vGFLRqN0wnPv87Y3sGOGtNcCwZG3tkw8Kae/XUgB0Ewd1t3LhEB1KEfBRvK
JPhIa+U+vbe8dHdQa7rx70Abm5v3l+TKoeaHI14nCpvX0+R6U6xYImsB4GT6ZMAx
6roPipHhCZEwaUZ6IFbNKBrriyJcLKa4FP4wjFS8oOImU4tFVM2eCO7vRyAyFMt9
ePv+N8GBMnqUQc5zl75wVEMJXSuvE0jwnRNEE0qZ6cTZoZCqqNGCz/UBzulcfn2Q
UEO6Js7i1AhHcU9piMLCFxh03QryktiuI7RoFFD6JyxT00cm17Z9CtGmE3fWBoQZ
iPrBFHmSQa8uu+HI0+Bc/E4q6lBxcS5+enUev8adAsoa8w4zksM3RO3zFOopHXNR
PChGR9uKmCD9qx/leYZ/4Fz0id+1YxYQxLSuQWYXdBC2CoAupzccfP8SdcepbPKd
Xkebg6n9CqdkKERpY8DXmeOSd1iIflTqOYAI5nWzP8mx7/nemLaNjkmMAuqGDqN3
RJU7VCymY0ogXEhtWw3WcYI6JSgnYbMBcYKuYJ1ktq70waUqVH8d1ocMNcnDInD9
c1IMT7V4mpQxHJ4NYCUTirD74Y9QB3fz7/AXoRRQOx8vBiAaP+Zwxtlrqz2V1qDM
Qzzc096gmb4YMKPS/yfuTiFE+mcDhtbl3uAO3wRm2Gs/M7oGQxRLp/uZxe+af+SB
zInSMIzFe6FI6LNEWusBrhDQjNBL/d1Tv9FYQshOg9M5IlGogfhOQFd4iDdUVpn6
7iMMAn1isYSCNUqMN7SLBzBnv6ZytGUUMWdoP8jNq/tnCquBrcqyXBvbHFIGrVyq
2VZOKjgPiyF3/g9Kg0FASM3kTGp7VVSTBpEOQgRTN+Lk/W/cse33opdlpqiypHR9
2u3XqFcbUDWVVRRgm+uumUu4HTjqyKEc5xsYDkgownVBSTaAWwlTdufsC6ywwpnD
pvmt/gDSLYaBusdjBfNrlpPyehdyiV2SNhWSGcmIhBQrRyrMjeDmCM1rkqQEthYe
Wp+7PhoxjKceYHOJo6vzu8dIASCezJdMjGanicKUzw+hYtflOiVY9ucw9sKyQsl4
+6L/XU19z7BrfrNfCjedk1LFbcgHNCzkEkIfoPLtE2Ua5dCAjpKXtp+ECCOHQS0t
zwIx9gUxr9MCqjvW5PfcpoGzfpi/LiEDUBWkRPoNnGH5HcBgiyMic4rxslM7B+nT

//pragma protect end_data_block
//pragma protect digest_block
lfIn+BD/XvLFDQ82V/7n9+AAIRU=
//pragma protect end_digest_block
//pragma protect end_protected
