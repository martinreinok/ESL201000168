// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H#*E42G!58YL\6>\V-54P)F;:8YN7GM5_"3\ZQ^Q^+<L^"\%(H3>IF@  
H45VZ:QE0_V+RI<O)^D1O)S]V,&LX8'._["/!#4$+3("X!#_OMIJ2'@  
H,5M@POL,)M4EV!\+@X-*R1+W2B"3C6I6V%Z^VO.._8!0(@EKW>^S @  
H+^PX.1$4AF\ U.!:)1(III )M_^\KN(]:"B5]<G:(S']FBNC$B&'G0  
H+BBKH%,JL>QW5FBN0@(L_R9SD1].B.0& X@F:V"&'RP#D?:9PA%JN   
`pragma protect encoding=(enctype="uuencode",bytes=13744       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@C#+U'&U_69.L(R]Y),:Y+_$K"6KQ05@IW!36&O+B=XT 
@4#R+8;S0<KL*GPESPIC=64W6FO%)C0'T03&*X1S\.V4 
@QUWOVKX)7Q>LNT(!&KS-)@O9^AQ@_K^=NX(_%0]%=<0 
@9MFP48FE@Z':HM8Z /.+5/+9("Z9$Y[>!*\73,3 HM\ 
@[1/M%09@K]6AJO./W\9^"^<KR:H$#9W^))U_"*H"Z#T 
@M 0.[A@3.XL&7VGA1#5[]$[8,C&2+UBW\=QF&:RJ9TT 
@3)7F4/2-[^WM^FI=&R?6CWHB]R_X ?AVNVU01G@Z'BL 
@408A,JNSEQ&8,L+!<W?![0*## BK2B"H.LZBDF7?B\P 
@O!'C;6%!L,D*&XRA*']?52;8\,>+!Y<AWYXO-V,RQ1  
@^54BB=4/U*1.54,J5%(2%#:H)HGU>UQ;,>E@0VB^DFD 
@*CN8+)90F>A7#A.4#Y)>>U[<!Y\>D&84@L,^OY&+B7, 
@](MY*.\-W15+*!4G1/F6&ESKZ(GD88'VETQFLCD"5+  
@!P!3)+4$:G0);^D.GK^6DZ?8_V0B(:SU6CFI3S='/=4 
@R.60)>7_)LY$+?4<E#%H%_I([)HTUHU?DA!3+ [ZFZT 
@]X8<?FPL[)(#!XF9>XBJ\>([W$O'.2-5Y*;^SA"Z?3P 
@9W#945>8!_9O[3CW 1'3O.*S>_FV@8H7D[';8@TO7YH 
@ G)Z?5 JQWQ$3R<3-=B1^OUE9S;5'Y1SR""GK,?;SW8 
@VE38G@YR(]M.D>GL(_R"N?#$GJC,_$#3K$*UM37TK:T 
@X_8T)EBWJ["J;<.$TB*AZ-B=R:9WM'$V@_Y3!:1R_-P 
@-^'RGQ"1CKQH0 = *BA3+)V"+CYUD[^0.:',*F^Y"-4 
@A?H;_?)4!M1!"@DG77E<*#5MG95JT=K$]H@UV'^I&BT 
@KOLYZ#-$$Q7\9Q3YJ36<.9,ZY&+ZN_(ZY #^8J>2-[, 
@38/V[/,#OLP15\""9,<3"!O=2AR/N<T,1T&.JT*#Y8  
@<\/[,,RR4._O+?0/0NORN(90OA1\1,*36Y[2E7=/.>H 
@0[V"_U3A^HLZ+P.*R'ZW <1=QZIV15W!Q%[G)48$6=0 
@YMDQ*3L/)P8GEL#MZU(X^Q&-C]8J_AL5(2$G,2OC\*D 
@%GNBN?!WQNZ3I$,Z<6^:F%(7F@$XAJ<:C/&72$TQ01  
@[OYEED]K$N?]MH*8$E]XKT/XEX%(,:1A715%RR/8FZ4 
@Y5WPC75<"[ U;R=TM2VKK&(%P+/):$C#UA?6]--JTN( 
@"$DB/^#-98BVB4%OIUNB0Q/LGG%OQ5HRR]MKW=*ZO?D 
@)Z<"L-H=Q(N6&TUT!"VY4];6-ZH R?NY+7D0I]+<*"$ 
@(?&'*GD>)?!MM+A$'EQ6_4[G>"%VR^RGM?TT+V"Z>/< 
@Y"!CBHT.K!?B.-BP+6PQW1:-...B4V,''<=$AS5SMW4 
@W\37#3;2^, 0H#?K TV_6?FXM#C(,$0C.J05ONC=OWD 
@ANF<6'QO%FR"0<X?4TF_X=AEQFGO[$_I#VNVDGC;W6H 
@B?8)%IH7U61PY-LZ*SM<Q=;WM%<K$TT<"=D%@JF$Z#D 
@K(HK.HK^C5>L[F&92%>VC)':TR8YCXS!Z"#3K;7PM1\ 
@SV@ '=D)>9T04GJ*Q^:L#$+D2PLA5ASD#+Y%>)=ZV8$ 
@0\3[PW"XA46"Q>_2C0=F>%*W$.08^S6QM0#]8)T$$#D 
@&P%?KG5WIU6:4>*3C_BC21*BVE"%NV.7?"?+[A58*90 
@8D#,"-HL'S6$A,X%_DAE*KDE#.L/(>UF@3"<R#_>BPT 
@3LTF^T8]<,Y0QN"P0:V1V!UWSO(DE"M09+HE)1<ARB  
@ F! ,;']8(LZ^5VN!=JSF=>I/>1P/!_X$0J-*I.0UZX 
@QMVBN<JR489NJ?TC$@IK1?;#8)_VW)PR'ONZ92R.H H 
@T@=PP^K9'S06/ZW+XY@F[B!:<R<WZ9$OE+[Q-@6J )@ 
@62=!<E,APC+2(T\BCHP4C<R2R8=PN0U0#>( 2/,?YA, 
@G/I<SQ#%F_2=A&T;JQB7GW $-BDT,J@QN C76J8N/O( 
@Y(10YK$/*';Z2.D*./ 6/1%2K+YJ-3U'/Q]'B$IK;^$ 
@E]X#(.96W\[_EHO,6;'9?NB*=GTYG]G<<FV/!+_KNX$ 
@7UU24JNWL <4<"U8P3,P/]&,SZ8O,U B\'>,=#UOKGT 
@257/3J#8_540IT$7_FVC^0@[3%*2'CMYK[J'J&I)E54 
@<X!WA=I$TVYPBLK\ICC>="%,@VDP$YZ3Z[VO0LXDQ1@ 
@(8/)2]\G4(R!\%-VQ3*-".?#02Q&9]3,YJ'MC+YT/#0 
@Y> YV<N'G,C.>)$KP%/?LCI03!LW;8XDK:V:Y]0Z$R\ 
@?\7+D%Q#Y:M*LZC"M!@Q^CMZ3 5 ]Z?'3HTOIE!X_*$ 
@D!"[[S6%]K1W=MF!#6-C^R%<N!LU/"&.$Q,^K4_MBL4 
@1B[2/J;BT9) 4=3%//R?%9_WG25B:!X(] J$?@#AGEX 
@@C@S,K13^MK2S@U!$^A@E_O$QQ&AIO,W$7^B!31 _,@ 
@KM=</F 5S8I-)/.W2[8;PCCO8AN _LJP;6&>R<:AY;< 
@-;L^+"DL;@Y@Q#&2\PE'[;;D?Z57/[5ZI)A7UTJO4HP 
@K?C([5IA\P>./?[-.1V:E;D>DNFEZ8P;Q$\=F"J7U\, 
@'1.<@F6+Y.I-]43!6W^ ?%/.*>(;?.Y_N*6C2W"0?^4 
@X!8#3;//K\ >]MXW#4W@D=.T<,LD(>_-_C#MZFGRN0\ 
@G",-9C)ED;=D4!1&P>^EQ\.Z:@/IB3?LY)RB*]KH L, 
@M5T&N.[?ZK_J+:;=<QIF.=:)L818[\)<!-_=4EDNV#0 
@,:K'J\-?&.E0P_8I19.G!A)0?4P7M>%F@/@O]_V,UQT 
@QMI>&8I8LG$ZH<2&I57YP.&N)\EJ[3$TO\NM&^4:"V4 
@/D#CRN_WZ"")PH%7K=GK@M.*C4X)LFQEG*N''=N=)Q  
@D\F)GQX3#D  \1&0I'05(6BBZ_7(.VHW')W'"=3'!3P 
@I?Z4_5!'^&WG#SF/J:P$KWIPS%^!C_VOZ@@81&_I>BX 
@8,61&"E.]&0^BC*K/V'Y@&LR)85 4+C4(97Q@8C5="$ 
@/Q1Q%0#MMMPXG@#U!,8(E2,LFQMUO9J^]*+NN"JQK#  
@?[LD2S#M]O"M*?OS=@A\H\IZWSY-,&:F&?:]YSM6'SH 
@KK2[WM2;?=.ONO!RECS1UW<$O&>XH0#;<%'<6YT7X4@ 
@' -[S;=30LX<$T2J!2_J$&<JF+V^+.RJN;Y[DCX26!< 
@EA/C,ZQGRV$I>&"# )D=RF7'4]^JN6@Q*I@(AC''DB$ 
@CWS)@1YVZ1M%=>"P]=I9$77&^0A.ST"9/I$W @FKDF4 
@"CD^!8TUV::!MAJW' KQ@9/=!1ZPJ;D' QL0<A:NAA, 
@\:K([P>B.M\.WL!1\H-K[Z*9(! DQ'[#*+DC:_?(.Z@ 
@;9SO> <AAG/(N!P3D1<")>JU;1SXHE#5@^3!/P>4]6X 
@0S+I>O/:.';B>!<0O2'YN1&2V^W'CG%I%Q836DZ+L8H 
@/'./-"+>) 6.;%1.K1LEWV_AU]]EO'9GU"<SA]A](!, 
@\1NC2R<\ZR2.2CJ12QDCXO1>VBB*Y0G8V-0UK>FIG@( 
@6)%;XJ 8&W\2ARRJ:OI2E9<3DSF$_F&^,]4C"F2&7Z4 
@>OY!0P(21XP>\HCD+98AA 4'>0U):&]_79-10YM)Q5L 
@Z:%G+$OS :2MYL;P<O^ RGH4T4NY9?=G*-G9MF<,@@T 
@\L/?4]V@?X$XI9?H ]_()RI4CUC$08]D#TV)KJDZ$0< 
@]C+4[B2+#\8 S-2L,-O#2@SH>LRN$7T-84?;%GXBBQH 
@9:\V')S=!MMHZ>%L?SJS+MTMC"X'OZ%P7IOTMZ8[P/4 
@JG[JR$1C9T7%#8!WI%-TLHYN)K- XB'HEI-E4R7C[-8 
@PZ3;Z0C<3[W9.-W_V\M5G+BIF3<KMQA O#4"6O:6B@L 
@12K(5<T'YY=1S2PU93+U<$8K9'07EY3QK+)4#?U@<_8 
@<TDEYF>8M$@'HMK,0P2<7I1I#IE+6I4B2J@6G]Z,'U, 
@<4TW9YH.;F1 /9*Z.,TA/E[@+%6B5F  \\$E$\DQIM0 
@;31*BK9253#H?7]F@L6W[<QU8$8%END@&"+G]BP$VTH 
@I%&EZ5.OJC"=QS] _N4J#TRFG2S-A>CWNIK^\,["FA$ 
@VIVNZ>WEU%:U=FN><;B(O@<"4W<J6JW025KO+DW5T[\ 
@&]\:!YOBKG%"J8U'K(W =QPL@?@-"R>!B -!UU(HH;T 
@%H7+<(%=E4YCM;5RJ8<92B#N3"..M.#Q/H6^J=MC,N0 
@_3J #';?_ ,WJBWU'5[Z9<:YE;O"S)MQ,\M,TF"&1QP 
@W[^P[&-A8_=6ER#Y:@W820T[3RZ#^G[+IJQ>+(FAIY$ 
@TR$7MI']F3/KO H_[2_8LF'C464/AS3:M_]0<N)[CM0 
@'_41KOAM:Z3BO>A8']WMG7Q3+<P@SP>=<=("(P5=4T0 
@*0LR\5ECD@K)@9FK& <S^VF\KLE/D%1/=6_&IQ"-M:@ 
@UDZ-SGTQ9A283$D R7N_$M&3Q?(7^ZRR7G8X\K.JD"8 
@U%[FOWWWN7"Q &0U:M2(TEKSIL1A"!""'0A1T5QLYF\ 
@RWYVM\T9HY<V$,L*\B].MD-]\QX7=M'KG\HR,Q!G?QL 
@\1PR=%FD_N*A.1'WS%*PVQU#P!.G&EG_Y.!UA@O-T'H 
@2?978X( "$X1S:M%7]C-&7W.Y4GT>;$AQ10I;*@>]^P 
@ KXFHFJ?9^MTY=-M:\?EH./U'K/^4;<;=/WN:9*RB04 
@)A3W[I%HL%LX&O9+?._PR0U-^<>*D%W=@U.LEQX(%98 
@@I#"[*8F'5;\+J-'I9,ICY(L^!4[HUN/?X3V3,SC61X 
@BY 6E6!O?VI$/8/07>(7=13QRNG"WM0*GNOY$RR'C!( 
@^IG,Q@R5.#$Y>W1KTB!3KKWANJ-_ )%J[;5<?J&JCGD 
@?(-K72SF=%;.R$GN.?5CJ\]5G*E^N.TX#&A^$OX?L64 
@?(^+,JNQ$.V=NB./RIQ6C' 2;%)LDT]J8!:C@UQQ_2D 
@A_*='LUY1HY[U,YAWQW06\WR>+9 W<!;)^NC=7)#PX, 
@GI?79=6NJ@/-KJ]_$$,F(M/1*U$MV%K5Y^>V@DB3'&$ 
@/RV6XO41C-UPXZSY&S*?E(_W2UC&=BU(9@5>S*X<OD$ 
@,T@+D^1?H^#S\T3.4U<<\50VP_Y]LDFUF/;!AY\(3*T 
@:+PS<+B(4 !9XSBHYY&;L/?^I:-2,[#$ZM$L/!;RRRH 
@EU)"6=STD3,V+?HR=COKYMD@:*:C0=64USW597=S7$\ 
@!QRC+?+ZBON+.5(I'@91*^':WDB$#>VQ?^$W'M/GX&@ 
@<'5L[BGJGV\5_ZX7HB)$!Q(W>?H'^69'K%HKY^6JZVD 
@8I6DM'SFWM[4\B':>7O')5_]0!ZJ0H;*7<@6Z7BT0R< 
@7^6L.Z.PGU\FU'[I0S=!.<5NSC[L!95K8=@^E-OO"%T 
@AK0-CHY:32=4V/]$C+>C/J=_WL+A] TJ! P/__3,BO$ 
@4R$*KT4# [#TF;(*(&3WA JVEY^DT@-MW0\A=:":4L( 
@J8IHW&AO7W7^_N'&MBWIF9!=2TUZ9+0>%6,<5HC(H^  
@NN3HPK]O^_[8D<J?W@*'MX2^)PV/)$%3IM/Q&8/EFN$ 
@84[LPWN>KJ&;#_,(<:2D(;:ZHZ3GAYL"WX<3TXT*X9$ 
@(2_%BSPC\\IQY$RI&3@CH:PF1;A-.?#,0&,<J5EJ&AX 
@B:Y_*R,TFH6UK/RVX/(I823B1F\C#I3N_J5F%V9)Y+< 
@H,;" R@7JA.?L-Z,/?B /QO*/S,0@FZ,H6I HG,_ DT 
@FD7?@::P^?6>*KY%YZ3D T04MKMMD120GB=#GMPBW)$ 
@NF[O6X"#5*"$ @!R%#L96%_1@<L^S1_\NSDYO_[F0:$ 
@T3B^GK_2-44JEL;>RK3%<%>0J.L'PS0=N):>E!4><LX 
@;G3(J5 2H\K&ATN)M "XB3_,?;9?9!M=,<1=K&_LD2X 
@2I/DI2<E/O94$:EBE%7TE,;ZWUAZ_Q&;F2$LYS4Q)=P 
@26?U6QL.KDWMU!)T)L]119-VD2\923])6.?NH-(7H:  
@-Y[":*8)CMC_@"6DQSHH4,0ZY=G\9(Q &Z<\VVI3W'< 
@R(Q;)T50.SLA3@:SIIR#9'NY!E39_ S55]W3IEY\"FP 
@5X?:Z<VV]^T(-Y+E\A2657ITD#K"HZO7G($D!3E5D;X 
@G^_%MJ)766[N/<\.@N58T2[YR0;+#!3)%_$S;CG7OR$ 
@;&/';):Y 9IM&$.SX+'<8NH":'/,'X#@F@X11>)Q M  
@YBX*@R*]'Q/B-H61UQ_K?$[^NTS*<TT69R:,,VD:9+P 
@[KZ5A-W' ;>$X]N]]&T:N_K$U+_-3G#K2:6A.EUL-D4 
@]1G:1A$6&KL[A8I!]\SQ6\\,T051TSQC@=R_NQ6Q^<$ 
@?0:'LK<3Q%OL8VQ[E.4)$@F;G*1K\X8_GIN.JEQ1?ZD 
@ZCU=8R+F,Y#%G"'06O\-X"@,BVX/=E+('"T9)^E#%D$ 
@7I<^ 70_4^2ZU9DR%'ZE_,9R=2?2;Z4U'_>4V5]RO6L 
@8.(U*B4@'Z'XF7@MGZ#*$5M#]?=%Z3D;+1ED+C!5#3$ 
@:^IA+$>\0XLZ*%*1#-TM6'B.M]?76 YCJ[+$.R2(F2D 
@",0H+KR'J%27B05<G?]F 4@Z[]SX/(.N/7]=3/]&E78 
@,J3""/@9YB([G.#S4W[)0<R.<<6DDO79G2&GJ9(L6^T 
@%7HW#V[]K T!(\<QGL> :>)"X.\=7,[BUTA:2,) W>L 
@!6*,1!.CF]>WH-)2.V\/9B@';E) :7/W+5$]X8ZZBCX 
@;?H;^! @H9894C44+0R:O\21^CNI;)X9>$)Y<=GAH2, 
@?KE=.MPB2B_=)R(:FMG>4]:&&0]/+$$I9X@3_M*4IP< 
@P3U]L?G?A&+?3* 465S$%@+?8#\2U7_5Y)GVV&JN]%0 
@VDL1%4&!LWZXE-"%*E:?(>-VRU-:5&PH.$L)D E%_6< 
@J0B1(4KA8L/A!RC:<BS0"D;M\:QM NU^EM#_RL_P\&  
@.ND+CAQ02?FH5I],@LL@05;>_@,)>><2VU)YN' $-TH 
@9R[!5I]!7/(3X.15:5<?!8 # 7@/R+K%(7"?=$A=AAL 
@!>/6]#IGD##7/1)VYXCK>T!;M06F'9;B1\;YZPB;6^D 
@,C-'/RD1]ZX P[<;<4&RJA#@&$>Z'\GI@_V4%X%P4U( 
@6'_'!ZF%,OKG/%&3&X,CJ4_41 >FC8\"ET8=O-.CU5$ 
@%J3V!$FK_ZJG<'P;5W3YAF7;$ RC@U8O*#/>2O$VCO8 
@UW#R?KY"%,[GH2-*Y/6.P8@T[%UF@S4UX>6,VB@0+"4 
@Z3#TMK]9L.1"4.T0P&\%N ;JX.A1T"RN.F]C6"%GU], 
@/.N3MA;E[SXI.X()4F9(N<9 )SR^5I?0 WC?4>9CU+  
@)ZBLZBOK6BT??X],66-9'6YF_?;M:2?0 O&<M/-DY'0 
@#%!Y+#;H'9JNFG0A&RU'!(>' HGDW#HT8G\P?]T1&-  
@%:KA-00\O":"?.T%=M&L5[GHX>PWHJR2 J5.M&W7.Z0 
@4?(BHRB]&?P+6-O Z%Y_VDKHY7V$AN;$%FFV4<&&0*D 
@YV^4$WUK-5@%G^!/]RN+N=O7O9:^$BVJW1ZF>+Z_N60 
@(4M@V3.#U= #QJRTX SF?M6F-$5?#J'9@>:['=1MROT 
@')5,33JM.@8^;5279MG'@KH@8R&FE">A.FS$FSK ,5P 
@39$W#Q>C($2TK\9+)Y'JYD:[P^(Q%V'T>IT<_BVA;L\ 
@2!63UK\FS6/OY%.M1#NKX15$?T;V6JB/9Y^9+*>%H^@ 
@MR:)EZE3S=T+:-RC:+\X?.LD+PW^5%F[?@2A*X]^U6T 
@B#?S[[A"KG>H,^M,$S4,&?$,%QYJ'# U6A]#7%>&-9D 
@<QA' +FWPP<?=-O2S"QQ8[H%P[J/[TN\%-X+0![][W@ 
@4-S%/:*1M[DJXS?-F<](X$-;GUM)VF^&8"-3K%*8\;$ 
@N^@YKO[I9( ,CDN"??20@',*TOQ+(2?I1M7"KSHH5'8 
@,[&S@WC "4A6 @:+[=7;H<"SD!(HS/3FI*1=2D$& OH 
@YJ/V:W!5E.''F,%37#/-?P2F7$8P/61:%S6J#6DIC4$ 
@OG]VL&VY3AQ/W K41,+F("AV?;LDRXT6[X@YH%"A23T 
@M$5R)NVG+TS?H/F^?+/^K3M+S8/,,WD/*R*L]'XY][$ 
@N7!,RY6U[KUL-=VXN!?U2(:D*-<9IJS'1G%GXB8L_QP 
@*#I21:E2S5%84Z-Z#-[8D3?3JJ.;&3=W22E?Q=P1]AL 
@%I.DE%NYVP08=D)<J2X]JY,0IOG";COAY<A*JWQ8O.0 
@_)4AE/%)\0<R0VIB^/YH>JBL5\D,.SN%HB3H?.I9+N< 
@5*2Y:ZOLI]$8I0(Q,DH3:S<GH2U?)TJK:/2"S!_*+WD 
@K5=J5R0W/EOF9>OH>2"475 \10U^2-QAF5EJ0&[L\8@ 
@K*Q2HA$9P./V[Q6WOY1.B#.8O4 ^Q<RA-GP(%Z4MM:( 
@5%_WNO$E-OUS#V'Q!-"YTI;=T9FAB$EG^ZM;9DXTO 4 
@.3D#G&FF]GO4T$\B=W)MUAH7$7)P3T2H/!9(M%4.U9X 
@\EM>2? 9)8:@,>(@PE9ZX4O]!Z46%V(S4E< .NAR -( 
@;L83/@AHSAZ[MC?R)^J,)H8?^)HCKB,Z-<%[?0JR@QH 
@"%(<PQEZK"Q'ON29.(Y$2@?=H<7!-A)=4V'F 7/-.2$ 
@LB4[/[F0@@%6:*K$@)8<9$9D.,OI@31$_:)D8Y+(,(4 
@>^ZGT!#D1H9M'WG8S K3A17] J%K\&YQ/7%XRS9BE(( 
@ XVJ3O\F4TN?#$7>P4"$H[)(<FA?H'B3)"+V62;O7!, 
@7TC2T/9$;R9^ON\/*C/S_*\Z*K2F9MO3HR+DKQ-ZZ3$ 
@2+EM1/'U>X*^6W)8/1I C\T/#RA= UB8H),'5Y $>7< 
@1;NZ5OA2L420LR18^OWA[AV@0T4[Z)E6E;7_O0)K.W\ 
@2VGV/6H?3Y9)/U *:[ONHS)4QH97(BL22YG@%2 X'64 
@Q-8X6,0W(00(*L]DE@S%$AJY\>X#$M'$N&)U']I_:%H 
@\;WRH'^ 'E:7_!^>]$*V.N@A$;:(X_3PGB_35?W[74D 
@3Q:Y>V='AQEU/SSJ$CNKR%BH#FHZJH_ MYI#4]TN& L 
@\S8P:E^]RBE-5C#%#U3'Y/^.3+4B\.V3TVJ:2&CV PT 
@P4BVNW8*IMKDBOOAX.3:LJ93?&,T"B8MNHJ&@[\H$U( 
@Y+:K\=9T,2#8RP6[5+K.,6Y ("OHG 6'X??;".<;I-@ 
@<4!#'%35+UIH2J/W=-%[?2$OKX& RW.Q.G0D_0D>:S8 
@3=#1*%S*%7\E7U;>HCW/["9F'M3<RX*4:G')61P-23H 
@H&A+0VQ:' @N!7R_/:W%LM^LIYXVA1P@:[O6M@:"[M, 
@QEX;L[8;B["2Q7H)YW"DVH%#28B9D3[.E%.AT(7[_JD 
@>0)-'QI4R]D-G&W!(VA=3P'N(BLZUR6,9!R5O'+J^P4 
@+M+Z.4UHNPKU4@"T]PVO.N5/J_H3O8_6(X?FAP"MJB4 
@ZE3DN]9-"* KB?L-YFK0"K+A4;T<D(B%QTQRET'-A9, 
@LM9D'9O[ZICE =D^(T^F3KF6/'Q3:<$'/Z*O]A1Q-&\ 
@/FG@F'"7EU+Q4 0)VQ*2):M'HJ9E+4*<?A'N<I(:5E$ 
@0^4_.&"D&ZGLA%?W!^3<FF=D]3+:A%%\V_3@<5G,&EH 
@@I>;]'@41'VFY!E_^7/7^1)/H.*D:"M7V&UI[D8F =, 
@+/TH98T+M)W\4KJ[4SYERMG!HY%\W;\J!,5:_#U5[2, 
@#V0*@=&<B:]GSU)L4^WB""YQ?G[\,B$%LDQFPQ2NL(X 
@ET*E3J_]F;,KSO):WQSN_S2_2MCFB-2^IJ+<[@;-,$@ 
@G]WO#^7+:"=:>+4X%CW>5(_"&#A3RI3^8C)W\U7>RJ$ 
@IE7\W\>%+09AEE/=;Y_*W4]SLO$HT&Z7;_EN@3V2WY@ 
@/2EUHOS[:G!&;5[TQ;ILF=T\_'PP->^HF!DWY POL\\ 
@ZUQ\KW FI@>7[TG&8RA'Q^1[;CWG(>XS-RB(W1 $N0P 
@$',T-[G)!_'T2I7DQ0GIDE/H/G\NE?/DIM'<!Q\P!R\ 
@^PJ',E4,NZ#IPGD6KV/FET77_O3&Q->4CX;@8C&1H,\ 
@\[>>7=X$ @>J2'DR5]?QDV12N[5]YW)ZGEO07-4W87\ 
@>Z!)O4 Y##@\K\TCB$SX$6D_A>3/@5.V'M.SA!?2I'( 
@+S?#S#Y[ST;/:U+B+6 #IY%.!DZ[=H);0"ICLNB:>CX 
@G[G@B4*Y!H$-G?TTT?W-Q@=A=3$K^EA^BD/M^F,V@'0 
@F:K(JH@'+&JO!.$QP%'Z3?DBP;7 ";SH'G]+R6>=\"  
@P)2"MCK..CM#Z)#[^^V"($/M;-Z906TA/65$ ''65 H 
@8<!8G7=3C=)@CJ>$=*)*ZT^8,E).43->$8/&")U&1\8 
@F?]K91I9(1DF"/1"KJMQ&G'^]TG2F?^!ES0=_'!;RNL 
@!F8OEN"C;MHR;I4]MB._&^\_<$#6U9/,6&"T;V\")A@ 
@WV'HL^R>H@YSWKN"'T:OUUGV%\ZMS=@'DXR6H.#57L  
@FGB=\$I]DGI386VZ9_@C.2:C.'S],12'"IF/@C:Z?*\ 
@,ZE*MS=OW&"Z/:9:"2S"%T$"(.SJCL^G7;D<\QLI*DL 
@ >9V&<3B8]-Z7@Y!DCD/NKPO?7Z)Q9U(X1^\B:JG80T 
@*Y#2OBY.I<1TM&]BD'7"%G'QD:,[4@.T6XS6O^?*R/( 
@?S=-]< ]%^\DE6.W70HIZ""ESD'6[JVRW>$?\UYD>Z0 
@[=?NK&&/ZVWO$EX/^-)UJG$#I%X1R<O-@ ZAFK[-?MT 
@C,*82W/GO$8#.GG5@I9XN_?//<DDA<VP^+L(C^'Q*"( 
@R!(ZA$D1#D$0B<Y!?[P7N0('NG3ZGE@4(3:BMNX:(+$ 
@VWWH)K!EE]3X->>MVGE7?X%P"I$[/B@!O=[CRMN9HRL 
@_ S9P*5^AR;EG?[C.QAK]<&!^JH1*C>/9KIJ4?)VXZ< 
@E<<QFW\^OK_:'SZ5@Q3KE>"J%LA)8QZD\P)>0[4TV:T 
@3/@TB2N6*>%*$ #$2T^JJ./EBR1._ASH+.1V_28-7]X 
@3_>U^8#?!+.:_&G],^NA\'V\?"$'!AFORX>'GL$]+ $ 
@S87$18_?R95A3&E1WL[V<6\%U]N>2'6D^><.+JYL(M  
@,QW.[.&BW'$R24GFD%<!HH*;=^4P?6]>R^MP7E=KL?D 
@D@6>UPP-SL!E_B21KP,[28D+M8#?D;L6"<@9G"F.T<X 
@\]WA)GN;K-RTE=JTT0LR1N>0^^TJN$&4AG7@1[=:LYD 
@!8@LY]%<&GG7Y/99_HM''VV6MYT #-).%.*/?O$[=/@ 
@7AG%22*'^?FSVYJ!8[RG?&7P]!M_L1H6R]H?PA/#G0X 
@F>=YOPN/PO\O^%2<8(0Y)^'ZQD3S'^8].'*6@8%"AE4 
@WZ;-<B*ZZ.EE[%9V1LVLO!;M1<JG3CK#[)H/N3T +<@ 
@43@)OIM051P8&[:0WB]ZSP^.V]EC\A"SZ#-!_S6\6R  
@K%3'_N%W*\]7:=1OV!Y_:<// %!(>\'USVTM&U!8OA( 
@J4%KHDUPT/IH"NUM_I%#*P/Y$Z@R59L9Q5_:XZ)]_D, 
@N5B.&8M:/C&9*LJP'V6Q^_TMY*>=&I3%DR%P-+COVH@ 
@3X$EC"\ZG4+1F;HX**DI657U)[PLY21Y?!GF06PI7V  
@*[F[2M4PA;#;@J;0B 4-S>1<-=QJ!5 )^B%B:5 ]^9X 
@N  5_ T4^CTZ3:EHY#('BM77=2JTX#KXU%R*AY0C]^4 
@B %32%4&#J 8I:53(;8,,,WTYKU+ ;.;Z,KF%,R\#Q< 
@+/RWI_G44->FX8J>Z2>2(BDM4LFQMV+BW;+N$PE2H2  
@O2W74<;:B*U48RS;S>"6BL? )KK4IE;.?#_*QEV7_#$ 
@!C9%\V]@NAMA/[]5"Z64*7_F)R2,/(JUZ/A:,18AWN8 
@L]8@7&;"#\;]P</.FIG- $.@XFV8M8MS61^FD_#6*U@ 
@= HI9,'O-MBC! 7G(65 6G2/ZIW*@IJ6[P7^Z#B]Z-X 
@GQ)$+I$=5R;M"4N?'3_PULY#VR$.02$B=5N9FLAEHO, 
@4?+Z[P:<OT,>&/P*(Q7YE:BK(TJ4YCN/.6A%":.V8C@ 
@*@*==&2YRK$O[,N07B2 [L:-NU4NW3AV1:*I!^VGF?, 
@]^6I0:SU%YJ'P06=T*7Y%"FD^X2-YRPCZ@!PZAZ&%#, 
@,4HP!Q'M7HW_(P5+L)L>'C=0 J:WYQQC7F7Q0E!.0O  
@XLQDI+X+9U.<7A2>O+JQ!S#.Q'I=GKMVRRQ&]@=?5WH 
@,PQ.>:]MGD(?<5F_$QJ?&QT5@YKI:SB<]43DY0^/&D  
@&5D2W& >E[+,1!AX%#34[\^BJL$&=&WP%8A-V0>E0N, 
@O"*<;XL5(5>\=,?J4$GBA  ] 7YE"MM]=-Q;R/M;>@0 
@6**O;GY^'S&5%W\$=0VA\%9<<QRY+;H*?:4-_;SDL:X 
@"F\/MMBF:4MY6^!<TBUSU6#KKA] X8'Q8K=HLXO-$[D 
@(03K6<2BP^QQI&NC07D=]O\F)83-_-D*WAYA6>Q0NWT 
@-@8J/'AEC[K-WIW+NRBF2.D-ZR4GFPRW%$)6$R\>IY\ 
@M558SNUZ/JDD3>W.U' )*#HU@0/J#(RI4LZ%/*FT-,8 
@<L=34^ -%##P<1+EA2>57,K5MU(A APNKZV./GX-=Y< 
@/_I$*E<,F%*6T,R5)P"-AFQN<T<$7KI6U7&Y5?Q/5#T 
@R:L^_E5L.X@C&II3;_&J^4 0)^(2X7[R?O]6+JVR/(< 
@2++:-"73(A,O!"3THC+-5&SDB#/,U'&R[SC^.]:J;,< 
@%6K<#->B&VJT1\'^.)@<^47W!<!5-G[4T@>KO.'ECF< 
@9J'TN1Y_X=E^%BS^'7_D\FI"U[ 4W@I7FN]V.)IJCYH 
@M;Y0+\6$C W!V4!KSU96B@#!' U<**RJ1"='<EPM%Y8 
@$Q%[?(1=(2.-J-0V)I+KS_^V8,6[>DK8]1U4!?F_"70 
@XE**(N'Y.:5 "LO8]U'8/X'Z5 ']7-^)<_&,QLY]POL 
@@AC$ _>+!7R@D7V.=8J>-S7S<MY!NZY>S<]^:!?NK @ 
@8NOJ)_Q%H ]XC:D Q_P>^1T&CFT<%('JD= _'E4^7L4 
@/83,$A')&"V&5"<B0IP4XP4118S)%!EY*7&KXHMPH+0 
@\XZ>WRUW/0X0?AYVGEZT[C=XQN4>LN5$VKL^9-;X9NP 
@$PK84'^=(VJ4120S2DY: A*533\"4&<6O=?I/HT[-'H 
@]B$=#.@B6!$SQL9$[JZI;FH&&)W[K0S.&_>$9:%G[[X 
@:TT/>2HYB&WMC:&K]_$@9'ZA$X=K.!$_@U8^.G##^Z, 
@Y"PPL72:JV(^+_ATCAR/>\(KL**<DUTDYS0O9<FN@^  
@RMK@LMKJ[->.Z@6"=#\=AL:/S#F\P4[)]$MMG2['4>T 
@Z,J6M?/51G[@F:H@2_=P=^<CIH>B>98,%C5-;Y$ QKT 
@\U>9$RT:&6K(7-2AI8!0-9?<%I-=DD%<Q6*<!ID85#8 
@$>(A3,H[0@/V$!F5I-/$T[$2,_Q'VS2K1/D [MRZ.;X 
@7L8[(KON/<M#$CD#34>8-KBV>4=8&5R(%DZ@87WF$\  
@V S"V!FE6\5C--):K5.&07&UI[!+.6-(#[[,Q@VVAFT 
@G8V+32;H0'XO$BLG?O#-K\0N[T\M/(XV+%A=9P%]MC$ 
@GAS7=JFCR!ZE:J:HAS9D!GSEVX)QS;)<O2\N_)="W5( 
@@HNP&F*M%Z6V6N!'1$F/RD_.D'V2W]<:P 4FJ;^#U)4 
@!85"+C_7&='.W32E?404U%1)HN'N":.[[6 ^?X7'#BL 
@T]R*?+SGB2&A>.EH:*:1Z])M< 1U)>25)8I?D%HKNRP 
@QN(M'R;#?NF#P88L0$VSW1L6HU9RCN))FM6"\TI/*CP 
@.YI$)HT6_[) )<RUSV'K.M( AQ/TB?3@1;A@HC_<X6H 
@^&C\1\\"<D-D_%GPU^(H;.K\1NR+3B:$8%ACP+P%XA< 
@Z"O>%S>S=6LYG?"5_D4# TYPDL._[:$>ADL_$7]3\;D 
@ %2<K@:ORG#!Z#T=:&?R:,&''>1(.U.80-J_3"^+J:, 
@9,N(ZX>5F57#])8.'/Q!ZF%H/27!T5*?@[I:I! RI*H 
@DF\*(#.]69J"2'PX5GN.@*>673E[;'1B'P,E0&O*JP< 
@ -S@Q#1+[6!\SJQK +R;RF$7_B]H%+B  6J%QYO35*4 
@H3]CC/;R,HQCP2.@%,U4<D3ORIW+9-S\E-S5LI?VR68 
@K:"R$(;3/%&1L)B@.49ZK -TWTN]H$/#^ [PE>JS'DD 
@<7;A5SVAR[J+%,F2L6@>2\-]%CB$ES-Z/&-_7)YG[PT 
@/82Y4=O>D02@P&"4"I.75/@3B=LBYW(K8Q7NJZ1S0VT 
@R5\9?JTK AVN3!L6P56D&D$XXNV^Q49E#2QTIW<K@YD 
@!@Z.TJ6L"D@&#S ZZS,V ,O#EQ^_7I?X@K7APS-C7%L 
@->_HP^=.S%S_L'?X\P$"MAMCLA[)S,A1%3ZB93AP[$L 
@#9C(P\B O')$0'JX9R&JK7ZHIM-E9AZ\*T;[AU,3'8$ 
@7$Y*HP*^J35X,3A&UL;;#)!EI=^Q'$>D:Y:=G1(_;S, 
@P)AN8/$[XV&6)&N<AP!C^*@5JV<&0P]M1D6NJ[[0?C\ 
@Q2G3!+=OZ9K[".1^Z[ M"Q+,="Q^A\LT>BK?7D\]KRL 
@+)?U?1(XK\)" &].P'%-RPOK^ZVH%/("Y+T8"H=!IM@ 
@9,_,3%RWFD'8=E/A^<X&UM+1=X6: X_[>[ %ILLH%[D 
@DS/[P *H;.V8=@BZ(Q!27SI$5 1E[@[G0-KJ++U..?4 
@Q5O]2K *USN\W.@/_@M9.^*\B/[]Y3\UGA\.E%@GEP< 
@TP+<;2&9/.'L"-=XX//>+ ,W]7R4^E%)V!3UWKLX.P@ 
@B<+<W3>T-@<KA%#5;;_B]3/:(%/K,@Z<*#K\;LE;PN  
@"18TF[V:V!2#1\X/9V9?=\=FX1C'OS*]C,OHCV1VGO< 
@_16[\H^Z1AH?G3R+.=?J4)ZZV53K)B8_3C.QN0OT<?$ 
@V_1!I3W"E1 ?A?Z#/6DJA&5[[SR1B(K&&O#-PCE[<B( 
@# H[2M$:^&)*9 \R>'.'WVU<MS4GFBZB(.$, *K0S4( 
@)6BJ9&3:Q*7S,5I#FRI1A[J]VYRE,LX[.)S/?6X"XC$ 
@I>3 $TRC[T4@FS.S?RFVDP^C3[65OC7ULK?F;U-=%B  
@#M%G6XC&KA@5]$MS<LP/;ZGI"R%,P@.JUT#A!?=/)6< 
@Z6<@Q< G_4/5H->SOAK["<)=OE^!#)=""[I"H-I^%(\ 
@@M#W ;V1?!AC0\,-G7&%G<8XW$6[6&QXF\H>CM*X3!4 
@%&G!UULSZ^7/$82)@:<J*@NL(S(Y'E!E=V5*,5QWT]$ 
@53<"<2&24=*I.3;VFO4W SNU]+\_?P9.6AB^1[/XVO$ 
@*"*3H1VGD;<BT1X7!@GEDMJPM@_,O7C0\Z%@>5@>^1P 
@F>+EI\:U/T'VF*0'3>"'$:WO]$(4%EQ(*9-^)B5)9U$ 
@!7A-O?S\]]<X$P^;KZ1II_09%FE/QBL7AVO%IM8!%YP 
@!OT\N %$#Y6@]#!1ZH1)_#<T%Q4'17NKC=#G:S3TM-  
@YLY)'9C3V43+/&IZ;&0^C2$(T,"E:LMU"L5K!G\6=YD 
@126[5R03&WPFA;RCN;1T_ME0G<F["7+%: .Q/[RPQA8 
@T)EX7>(KI#23(\$F4*L"C#=E%7I[M*TL.2\B;:HYC.  
@O);0- PR%+\7^W!ASAVGH3$(1IQY7FF=R*.O]_5_FF< 
@JS_6@-K4!19'CEAB#6=ITRY*+]TG$/5TG"!:GL'S[<$ 
@F LN,AHK;^,D85_R=;IF@2M7=.BJUA]S%POT.@5%P-@ 
@32QO(1S,6'_VB/]VL 1Y1K52B0@L94:S<05@PM5X1_L 
@GY2%\1AQL?XKA1 2L30]L27KSGC-51/V1UP[ /YJV!T 
@" S&H'F*]XVW 5?V*K:QXQ//U;52+?F<<ZGT^,NP!6$ 
@4WJ49E-;O3@C)\4,U/I7Y2>M5:UE6-66:"IBL:_J@<( 
@7O8+*=*YGKW]%(VGP#BU:9Z@]OZB+]?&TO.]"/QOM%@ 
@^V_5Q7<^ZEK/XG^:)Z[G/:8F/D=+A[W!V:M.*# +E@L 
@8^?]6?P+T[TJM@TXB3DDN>+0-6S]-[NE&%_C*S^L6Q  
@^9T.^L1N*N#.=L@C;39?&;<<5R>5/31<&5G =)IUS]$ 
@C(3'0> SU!W]X)3BGRYU,;%O1NVL*A"FLAK7%DHI>+P 
@%52L^!<&K+1U%1KM\)?W\.-G-!1S%=?E0,0@,DU;IF( 
@)&T/0S>+#@Q2($'6)SX5H@T'%7JQVZA:9#@U\&5:7@@ 
@]Y'6UGD^4&I0#!2A55 /(-^5XPB>!HUUNF&&8LVM=[< 
@94'G%3QQE$QW7M.3_YPRN++I"AIWS- P5('A3Z4 MS$ 
@PA=TQT]<UE:ERUB]D!)F92**P?H:4V9D*M;VVC[!IFH 
@*0<GV".W0+6T':[[O_&I(6HAAG^MB4T+>_<Y-PR2_.4 
@YNB<&#28FM#4SRU!72E,_/.&&,Q+#TYR0-NV>!RG7"< 
@\7L*/_(<4'%&Q6LMM0,7.YW1^,4<9W>Z.J5_LMB?HY8 
@$@/9T]OZ-R=;1C*F>%[1GU(G,II@5[UH$;$XO$#%G5X 
@EI0S.K]9^.XVY$S,Q35W[RB=WFETP4QG\%O>A]8S%Z8 
@_O[YS,Q4^(;Q+/9RY&MQFZDI$9S5:)>T!P,(=;+K-%$ 
@#F&1G&.NQ,26AT36-+>=M$W P@CGV+BZ322#G([U,3X 
@%2B;A#XX^FJ=;O1[BHXZ/:'@=$#*M)+-N(#] 7!87V@ 
@H?>MH,:VVD*B:>94\T-,$XX>]C:(G1H\;@2U*55&+OL 
@MT&Q*M- !BE!FS1?I!IO)Q$\OOAIBSBZY\X1RI81Y98 
@@+:&RFTK<8H4-NG<L3DWC+<1]A5[SM8-KZQL-X8,C/, 
@/)6-\U\/ &I[%)[,%'*'_AQ3ER"U2M'G-'_NQ[MIZ,( 
@X&%9V <1\*:K4PQT;*VE?CW(V%MQT]-]70\T*</-:/$ 
@"CSRT7E#R8-#8 8'<8-0'<49H"S($A*L_X) ^?ZT'<L 
@KE6O?M5V&D)V[&7OPL6=Y \HA4L ;3@R8=13!,\:>7L 
@L8G4)ZP2,?=Z'1\&UP5RY?/G%1;J(*,<#._,__/$L"< 
@SEN[&O>H$BQ_45QZ@D6(X*5CW*YU_T8(F%UNS>+2"7$ 
@ZU;_66!JNDJ^P\.^1K%A;Z/E,5BAK)P\D'"$A-D>]=D 
@K\ORS[%;[J;R92L_EM?0U5,GSCH2\/X4(G)4;F3D5;  
@B%:O@T+#Z<^W"Q17K.@QL/E9G!$PB<\=@5HJJ#VD;TH 
@5@!H^JZ#Y%2KXT&K0-]3M"<<F-8%K$P--%^N^*VW("0 
@\)A SD!,7IA,_(0EKD%4 0C&)PX?TB%1;\Q#7L7+4M@ 
@W:K.N'9U9JPZ]+G7[42_6M4GA_@A\H#75R/4([Y&#U\ 
@T@OF#NVBWU4+^W"%+98N!R=TQ;NS[-3G.'P'D?0KJLX 
@7K.#^^\= Y^0#?M_DS4>1,ZGV;5CIXBT&:?X'SVCWI$ 
@7]:!\K3J8(KY1_M= XM \T!1SBS:+@*P-$--,R1^10  
@O>9<800P<7R-< N\E=&%>N;P!!)+\\C2NE]>YB"7D2D 
@;MV.J25T\X_K[8\1):&SS5<JDTFP_Q.8I]OY0G'$</< 
@S&_A""$R3)*IQ*E .,:(F'\ZI4Q4E5NR%9B]XA:<M^\ 
@"@F!/[=\1J$-?7JBD(<\JZ*FV(G!6J]D4ZVR%M7$^D8 
@;;9\/ 4GFMG39+(9"EF[&FRF-L(:X4^J=*F0I<U(!K, 
@WUJ8QR,I)QTZ%X(=")VR00._NQY]5@)RK F13[W;&Y  
@=FTO%[<RZ"VK/=<M3]Z80#-(Q1=[0]K ":4!R583'[\ 
@!8I?/A.8-[&:M9+_"*D7G02TZ7QDU0LJD9@L1PZ!^^( 
@TEN_4^$R=)\W4V\XZDJ*_Z2&;(_J,&3+_VJ*,C2D( 0 
@LJ5(.:A2'AOV,2"[&'\_'IX5!'5/MV8'U2D[0=/6W , 
@ X?D;KA!V6UB&7.9TE;XIOUR4;Q5/F8<0X*U_&5!NO8 
@,@A<_$2MPMXW&?X />H$+L8W905*V_'U^*LC0??RO38 
@+ $RX'Y"OWPAH!8H5#SHE8:?BJ .YXST:1CVKW&<+DP 
@ 0A3D]9A]4(,R55(1C$[2V&UJZTR0!V!>%H/3['>+LD 
@;UD2I=6.^Q8BS2 _7#N8:ILM8 :Y6;E-]VNP=LI#M7D 
@6:+>(48&&S6HX%;C723!IB;E"/%Z[P4I![B]&K>(GJP 
@5#IS-UU@]SJP'VU(!_G(-B-G\)S(M$^ +5S:$Y!%C6, 
@3>B9'8:L$Z1[HE9UG>ZN1'95OYRGB1W%HZZ9!:Y0V!\ 
@RR6H:^% D P)IUWIQ3%,>0>0 M+1-@BP. /SAE4/K.8 
@WKTW$97KP#)[5UG7S4]!]9E4YW03J_0[>,J24)6 MS  
@;LO$(]O31=^&\-\U49T?/VNE[\*VTL.T0.5;:^G)Y1, 
@ X!OU_EMZ+-(22F(3W.M'IW6ZO&19;-P)&>)G'-O:H( 
@M0*JA@!)6[>U<X1?7&*I$G-AYV533P/+V_HRV/IT_7( 
0T#'QV#=MJM,WJM"E+;_RCP  
`pragma protect end_protected
