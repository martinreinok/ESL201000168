// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 03:52:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eISHNLKlVhKjKW+rl0FiM9z0PJFTfRxaew3ajDAuDa1wIOgULZ83wZ+hV4DkEAmJ
HMSUNdUf98uOWnO4hcM0CLZHBsQDZVlfd6tJHYj+BX/zJXUPkuUYc3QvgdGKeirH
tK6vXZGHdObeUpQ463Z+wCYwGj0R8RyluQU2Ky9hejM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12656)
z744UsSOi3dSsXK9532oEtcbs4pqdUSCPurbvuQPJQd783qxr10Dy0oWyVbSouDd
NbkQauzM4Fxk6epLbLTqVLTCPGQummbaqhnE9fyqZPUl1AIYFCY71W0E7mBClDCa
d3o5vK4HLykLpQCLEpaLJP0QcuAw5iHm1BD6cRViQxYL3OY39DsTGFyE6Fpmsn9+
m+rltfF8lqeUWnjHV4NSz36ClrPnn9LMOBQ4rVLdbYWLSoRtqOvWYHcYEPkYfXlb
RkI5Be5ZzzhaYyhB+za0e1GwgVJqfpXVmnlLts8EDJFZOt7vE6HjjmPO+CAVNILo
yEeip9vwrOd/Ax5gAHTXSkk2wUMHQWyeCMW2lA+iaYUvOuSm6Mdqq8UdNtL4cdnH
tCeKPUPsOUFeACVR9lC5Zj4IZusCd3TF1Kq89dBb3XEGKgiFdnSZwx/bqt13ght4
Aj1oR2KTAmgk3qRkUsq8hFf/LYf4vQ8MICVC9hyU9CrN704yuS2P3fo6tI3VOIgK
NU8fd+EcNSnIr2JqnPDdBExcsxuxL5PKHp0NEmuTDoz4ofo2/jfZVutaylFZ1WDd
HIcWmZMoCPMr60pE98b7AwMMqTsWoWSZfUXky3hSlV+uLS33V4R2Kr6/JU6wi5kc
ltYQh+zSYs2aNscGGP4qDzlHcFEKtCGQpZeNoNpJ1pDho/0KvLPR+zpVFOvSUKw4
jHdy49xkjlyvcGW2t5q7sEKvUJG2lPOYdssNaz6+l1msJB485EZLt7QRh6kFwvc8
g+WYq4vXeM21wLRDDsgVRJQSVas0gcBQlDx8t8+mHhE8X0e7z7oVGUWXmOqPCBlO
2xDcPFhOM3qpgHvnynRfoS9KdtKEnT3/aK3Zo/n8uNEU6R7Zmhp3/Ao3mwGfnz2s
RNFyWHN2RQFfp5kTxNNVg3Mk9e5+Zt7vR+TAXETrnQqLwGXWOCMvxpQHi5da1OqX
dXBuD5lth0Llr94EUjMi9/KNcW2OuCzlUOJwFb4ewqjG1CDXxYdIkwgUENKGaUTt
lHoXylUkkcxXLBz8UbZFlMCHWyEuor0f6JDjn3sCYXnBGmGr4O/9zcaQZGyquPA+
/FAJyqOSnPycEjsooHGdkT8Ryjh7bC1TzcFzVfYmOrlfRZplHxHEFXM1gpKwqx+n
7hTTRfY/lvb/clc0oTVNuxXd9t8QSeXRaARhzgsVbIcflhGOj6z1o+5gHHjUuqbu
GQeSroXBLGoLMh9Vd+qzMgwe8lo01DDmqLaR1j6UH0dd4//0Sh6/mdztKWFvq4jS
b7oeHlamcaixvk7hYj9rr0lov33TpPFDEQNms2HvS/d9f/j+aFD1ZgrQyCNNR8qj
hv2BReQs/3YmMlbyIgdewMj4iVaVb87VHKr7S+yXZL88HPa6Nt3qfmy92MIoZbIP
eyalxI8gHR7hDYPx/EkgswhdY+DvGg/rRy3R5qkp5UccdTQXz+q7QahG/t0wn4gc
JyFdpcufshFlM7KSyaU7uLe5vZvN2kXfxz/D99lwxZKj96a6iGXVZNXfSc2NdBb0
Zi3jmKVFmqJ2Kc1N/ckvdEAmfcr2SS5ev7pMur9PBEhVx4W2lc52SDvGcR8BG175
8Abt1EnA6rC8qzHGl9pU40FJ9kg717t66ll4dL/F8Yi0pG5LiZXuo63BQi1tzSBs
PEiUQEdfMCK7jIPEqqCZJn2BpDZ7JYSj4F0DgO9kNTsKRmt9db2e6gg9MAlxme51
fAZyPZnoEqe0Df59xdvUjNEFDSuBPDOVDDSs0p39VYyr1kiSSHFIfRIf9HUGdL+J
FZdpZ+FFObi0k+NkzqnWLSWHQSoIsPRey6iQ2hyIHr+lztagzaKhxWnUu10s1FdS
FtzdBTHSVDQ2DHRo/G3MEgYOk9i5gQ4Ub47h7qTbTaMILRt+T2hZH65L8onSzQIm
6GTu1303e5MFnLsJ2aFXOKBm3cuSOnFe/WTOJXshB4lNtG910Iu/eF5rJg0YvScX
MikGypS60f/M3UsLAPoRM+GYp0EZUMfjZralGiNIOg7xjSo1gAldfQNfiZXG8VKL
m0d4UCEfYpoeFlnDAsocXsGJtb6sBdUKjQ089BvBaHICEwP5A95DYTXdMmEceROf
0ha/PK2KKCeD2AbIvOOAKQoyv4NHugmfyQdONAJj1+Op83KLsbrLU/fF11CcPKBG
CqTCGKRaZtm9daF8uCyrH5F96rzrFQucIRB3JMC6Bg4Pc7fmNee3KqKcLaNmZmQw
bInYd9sA9WUzmq4/Zw42eDWEyJA5gfLxsj8KpNTEcifJ5Fa2Py5lz9619w1u9Cpu
P+4ws0Y0fxuKAbs9lsIp8Jb0zqs5EDmkRamjOMbF5Gjg+0kpVXMyykVHH/GoVjaW
kdhauEYUYOrKCNX/m9tLB32sKcO/InYLvXhQYwkXFSG7kHIm/E3IG5aYPyi4Acry
lA/lyhQMQMhcMU+/q5kzwT1FKEZd17V41BM6hTXBzrdFWbZJvyGcWd4CLzLRkozD
YJ62d9jweNwQlp+quQjRsUFDJ3kAGgEaarzlscImqAP6TBAS0ORtzZbiVq9shJw+
zaswCnMG+Hb7FItAK6EVdRhcMgcF9HVz67iL/JCiSJJMx8yeHvISDeb/1j5axN2a
zxyohnMQ2YgVh/h3jxZmebCBb6Rfb3F/wD8O3t0dzUfMvFvHP/c/12Y+Qhv8/VXi
W4juhFf04nyL6M9+X6MSKliuWQznnTFGKBW0wSPs4uvLTAbGfW3cBbFwTWq0j/gO
OcSe/F7hUjId9tEplnxNijyInmtFI5qogDA0BK3wlPxOp+iNRUPn5xgUr0aiG5Dy
G4naFjxkGllPtBAtdH3PzK67SDrhhBS6oKlN3EzcJog4MPyIPjVxXLSDmbqz6cZ8
Vzx9Q9gocAp2f8q25X11wrypv+l/dmrpujOFDbDfOwG+ZXNT1Pr3ooNgvKqhBVs0
u55wMtfqD/iE11gV7LMNhF9686ptwqhm2xaGd1g6W0JMb2a109TeC3r+ypt9OeL/
Qa9t1ZRVHchlS29ltNoBXQgHcGIhDzcDnvkiUoYbRrsw7xnz9plQgOP0sBQukU4O
Mr9fH5YKInzVpJgfvUmLJ4nwhlNS6M4Cz0d8OVLFxsTHzxAnlNDchT6Y7Or706nE
poTouyzjBYiax7zPSPD6OcJllVvyV4uGjhDhmRx7iN9Xj8gYqUsG/Vpc+tZ8Pj7b
2e7+DiPr0Sy3eSFCqIpGPBmnu9aVHtVyuuZpLHxCJt6STkKwMDwSz8G0dXW4XGtS
evLemeFC0kMW34uR5GbK6YFhUJDZrCCK5p/3FRYOhoXjebr39INw8ek3xcNV97sD
o6ejw4pyVdrHy0zdLh9q2EETfzWRxqux4f7WmvfTsRdRK2WMIFZg1WePnq36PH3n
s+BefSHD0F/JskLJstcecldIY7xWCIrlsvVaqafRTq4bT05xS5OSGEs9++qHsXV0
iMomkIhfobDsCLNuJAj6LBF9T09p4rw7Sh5FoPqr+KLrD4uhIWl5aKFJ+LNnjr47
wzDIIWzc05KB3wOAvGAZ4yzQKlQgN7F41tGMMhpySIEME9CDmeCMjCA21tdzbAc2
dm/t93ra6kz560T/0IDQwdV1YfglwZ1CW18SyVXBTdsz5OSrampo2+ZCAc31WrMP
4rwBFpkviMsq6gIQe8XehM/pVQEiq90j/A6FjheOk851IC17CtGJpyVL/MIdev4N
n9Zd5sBGq3RoGmGUxBE6q2jtc/86satzAyLfq1Hq0TkZ6WG4d10r2ct+7iysnafr
hWydo6RCpTJAyYzvaHjNXMK+IypbnPQZjse3b/2PGVw/5YZNdoF7zaPJaJygCKr6
T8aL6OAnUC3QsyuMh5m7iOAv3BJ8YhdJhnp+2S5UBaL4bzMfNjU0Hc6MR6glTbpA
0IZV7W8Q5FpEKvDVrcSW/A3ncA/Y4mJIFyMeUdP31v4/++7pStjdI6UI9r5eKmNk
E91wyn6uD1bp0G1CTo6YwxxHlhp7Xz6eqvRCwwXnYJBxjmnTxTTaz2rclhpjVKIm
jXjj5Cj/gV8yEzzDmVkxExLtnp4jc5h8aSbGCByY1LtryDiIEeSvJbmWEvWyeBXw
YcBAodMuBMM3SgULtrQT7C8nvYToF2Y7W7CDqL3/OnCDUSKAFcVcGht1EcDeDjit
zLNBzvhKfnX3fLIycnF1DmxtX0Q2Rm5C9IdIZnzBD+S2QAPYCZ0TQbWyM8eIzNz9
VG130d0FrgszN9lnqf001FFJxPj7tZX+YfmQNXJ9GWvAL8FOASK1W5hzcEQUreMD
tlPPRPISFTbv8m+jvExzU8eJF0zAFTncwwXRF+essBYA/wfX5eGKJoqZRRwTdXES
jPUNbaiXh2IWSjb7XeYKOgknekgyC8r036ni8X6+Or8mXLLUBZqIBCow2gRKXgq8
Hdg1cYe6fUt51EyB1bVaxnAPCJjLMpBjTbaKRPQxhR4v9lZEzVIezGFwgdJVkJev
dU/s0mcishLGB+WMe5xxrDWarQThsgCt41+OmTlYLvNBBxbdwUfo7+PWUD+0bkSB
2k6CKkMBa3+DpiLvPGBgh3t0qCcYsu+bVIBZIajixs2fR4+sL6dXl7yHiC46J/aF
7WLyAXeKaLWwwNzICcQmydGcqmxkjB53J06xhfGiji5B4aCESS2t8PTnno9jKGgj
wJUFFrVslnXdtQsfs1Hju8UBad+prRuKOc2tEREicxEPoObwXuMcT6QqVyUzASXU
D0TaAKlGfTsp/Nl0O4O0T8pMg/58v4uaMTX3ifBl73HD4BRLn2D9iP3szpYPG839
SudNrN22Ok/QaGAyTVuPAVp6FICAQy8tU3c782FjcQmPdo2UO9VokGyqMmm0lO64
1TNno8TxzI+NRsKdCZbyNf+V8qD8+xkiF+6BNsj+xf4piCW6PHgDpEFYRlTtiteZ
bV110XRGM1eDZctUscU052dNGLo1GYalCb7VJQtOkrF4I/ndVWm4OoxBP5KV1m3+
X+T+aRQ4NbqrCfJxuXJavvCljAQjjEcOuO6wVoLzfLHDISOPTKYO6O/gymD4E3+M
itkf23xd/eAK9t8mbw9lgdxEttf/a4tGB6ltnuDhlk6V5eCxg3MXL4RHhqF0N1ut
RDgGamAoZmgKDAEFSitJld3bbCJFJ6yLVofC08hSb8fnYEofUZFRqqvUdHzVxcWI
x9qqd5OULK3IKUG6GJh7kMMrz8TpZ/elP6xgUtLkUa1tpLpH4gqBqpbexwKeEYpZ
sEiNN9DMmDtKhmev4It2tqc1pvqvOAiAXLUGbfReBrc/EdgUk/VSelyo0sjq1OXx
lp51bbC9HEdTJmBWvMQEwopeyB5LuUBgbcmv+VbqvHzAT4vLzOZgcgx9mCuscoDg
RxmhBtGrhTNXDWhwCktgjtOJ7o/7W4VcQDnTytwO9XmNE3xCM0Ekk4t5DFD0+4Gq
uu3RwBFO16pGoXYpyaaiAea9sHPPRdya08sR5yuGCReQYfjaAzrO7oA+FHdpgUi5
B14RIa492g0SMCSUIM1xY+bKdVIS9FvQkStR+zkIG5tVs4w8DghgBTvFFmwyrXA2
DovszhwNbU74Wqc7gfol3pwf4UuJ8jbH+9Hmo0JpHilOLLRsmXfcjiSyWBV/Mrwo
ZT9pd8C/Xam/AqtayVawQLns/uBJZnKcLpUp1OQ+VoQO+U4pB1qLZ+1P5UzLdMeM
d2pstcrFM6DFee6gYVCSyWaG7bt+RAww/fmKgcNTgnWLrrSXWqL4tdiACwOY2A+s
k9uzg1blqRjF2+uy2Lb3kj1wY3pcPx/xHRoUoQPnxGZvAuoUVpTDl5mbowMFqCZ1
4oHfkObNcBnF1YuAOk036h4NmK1Vq0gQyPWmrLHLrwh0hgY1xMMvCfCSQxgnCHpo
egCWNhyiw1LXxoXi1sF/7Ng5DBgQ6lXAFOWi+uV+udQS289EAYdkM8va21/Ska6j
rxI8AKblEqi6faW+vAYc1VgAYZag22iaRFVEIKkxz3AYKgHAE7VfFGfieA2jblEG
KaV5ra9G50xB0Yjs2rmrryx2wFGUHbczGKqZoW3JrcID7gKEH4KJ/sOBs9laSdTd
Gge8o4uslNfd5eP9Lw4nhWi90mMgGwVaA2WuBtN6zvt0+PYzWLpLy5nd4ii91Lbc
REL52UB94atVcoIaNM8qwu6JK7ZWt9yQvViv27gOgb3acmBnokK+2yzvievUVOY3
pVPjSsaQKHk4mZVIyrdztwwh2gG+whHp+L/RVbDl8b1vCMz8VBFYD5YXVta3wi5V
h/kzsYBB3I26JNoh4OURXoBC+ChWTC5STSgqDqGnd3j1xmqRZ3G+e5CYYXYV6ko9
NuQUbq5zMYFLeKZlFZ8oq08BlqrwcC4zA79AtjnFTfMWM/XjjMUTxDL6ly75LRYR
qzKCqmez83HlhigT6C1y3Ow1rhREpxfrN0PJGL2fkpU731TWPCItE9pZERjIXM4H
LDT0qDU0kTk3HAPoJA/0Nl7zNjhx7X3bEkw/XWH2uAUxz6VYwOCrKVzRGImM+BdI
sLEjgbOZeTl0YRK2MMcLA6uFLYqhOEVpVgVl5XimWHfObCEAc6fQTJ66B9IrHsED
uoyDf/0fiNV/vq01Xztp0wuy7/G8+dakrcLsRpwUwID94HxOlMDnN811rZBkjeos
Z9AkJR20/WBDtLl7tW8h0MEXqyJUWfANYwUxRAltjm6vYy86ctG3zXsGTzS8euFX
rXx/zMrbogCefPzc0C3wSlXHZgpwdG5e3gDEYl0iSkRsIbi9trnSEYXHCFvp83G1
ZEd6XHLt8wivIK4u1pMbp8ENE3btgYKIRxvNuHCpkDZhjhRMrsDpQXnz9gVAVxQV
vntJOPKpvNhJPOosWDRxnDmdFJS3xbXdOmySYHCwAHQKQDJapdwo8QnMnP8dw9w+
N+Evq1pLwcMuG4wRp2gKfkesXlilEcsHuLuXXvmYM1qiB2ZQnhEk9bFYXnw+s/sy
3c7gf3ghVkkReUs4AJU8ZML3BuCXhLzpe7/sogdHnCCmhEOUm4QA9y0Xc1abXKPh
HKl/cWRXvJJt+hxbrGFWKlamdWaDDZgAUIslvq7yCgpgRHXsSutVYqJQFpH/s1T4
iu51H08YpHuHJCeHgky3Xy8tUIQGjPEMISn7lE5BH7f1o4Rxy3Jo9i8UpK72pGqp
yyi3jc1D9ymI/VIpHF5k5NJp6pRmogcctI1n6rrDlhNb/isPZ6ReXo4eMp/2GOF6
1TnIIhzTcQs6VlPl+IiEYZmAb1/7Ql2t35oe3vqYnVc+Kd3QEorC4GQgLkXrLBYN
bQh1n2PZVYC3J+bIxyZlt/P01XLFWV6PyrSBUz9Xy7dqEQnTUhVHq5Jv9ySpp6LG
l/PsiECu3C9tzw1k4+NXdRNukVi/OnhU1+AL+wSfv+5quQIsK6TZLTd4to1NkqIK
8DHCHSUoL8Njvzo7oZUnsHRYqRtHRaZiJU65L/GoFIgk4oMl9Reh0dN+tgRvGV4f
lh5hFUxDboEesmrZmy+s+gEycpxBBO61lwEqvwRbpwaf2zQnrt96knmE9q3ro0l4
ob33Azlehu/SJjcXgNmV2f8dSmhxtEtFIw56d5YQLNYahwxJYeSMRlrjb4jnbz0a
2toBq/0Zajrp+GhHVoVIYwsNzXINIjMCRoVT5dgghEbwSY3GRl/K7aLRC3Ub1lLN
mxvSg8J8hiNgw0CrYzN5izE6NXWeTXyNY373v4eqRw37Bz4Dh1N5mXZxDpIMJGJ6
Qwu7zwYLAq04N1ig0op3iikY+0v7OeqHEhKlX7lZFMGevf1pG8qt8ksd/c+sa+Uk
FgxAJJMLfv2pK1ybr4VpT33qW6wkDJzxoJ5NIN2O+rN7JGQbLFcJaXxcXOmWrItr
dTENCt9FApPSiM9PIKsYXBh52ey4EM/LvEyYe6o7rw63fImSXPCehhuIzp4MGdaL
D6XcHOyLwfsudWGIhd8i+BW0SGYkPnw48W3pt4ug1ZztHTAxhzoUbA6tlsu8HIFK
uOYZqCuMVYfzu64CHMAbivOLoWrN0Xu4GTb7THCYDoDgjKjMrAwPtQXfkZs6Fb4u
qZP4wiLu4EvpQYURiY7mvA9Fe/BEjngh8oF0e3+fiDsELFjT73MU2Zaem5mJsJGh
lDrUbgDFZypHDD1O+TUNrPEP7SRqC1sAlAkELF3D7qveJvMATsu1WE+gcXjX32Fu
h/c5Bc2Swz9/wg0bl17yphE6SIeuUhjWGezFi4Uc2qNhQaRHmN40carsHpreooJJ
9ApNxat23wjN+xJ9l2hVjNk2ajaggNmsGMW0cPjcfw+aybMLGUAVPHfIHc9yN4cn
4/umoECCP3Rkitl/u+5MIqM/Ybwjf9eSpmBkj8LUpW0Tj64c7pdIFA7fLx1nUF1t
uiKSylu37HdJWZxvgC8BlGlPkDC3Oqn1cql+7cnK6LUrEJewsO0ZB91OVv0Tr9B+
DZSJUzCfRl1BAuDTIrvOIoAu45XvrK0t5n4md13KJ0OrVXsq9b/WrnBIoj5Hz33T
P+G5HdppdTZnxeFXfAyM6OZjuYtkDbg4WYoGXKermQTdnEzfDLjwFEEMk3f1f6A1
etHKIy6RJUxrppJxTCCF2hmb15PY63doOzaAntZ66HiwSauhYrhG4XWW/UBMYzkm
eX6v9fzBRlZ1iTXV8nGlOxEE08FmgDmXg2aWlCDYSiG/qA8WCjRPut7r3bveNsjP
N5MSND539wjocq77SBHvF58SxMMBqIrsC6NocqGkJf9F5BtAexE5BzYZcAgGaNHN
LukK1xfFmPTp5PW92MNbfG+ypO88ga6EIjxss3iseDZHx6DLDm0UXytLbFhlw0CU
HXK5UvGUr161jcFR8KwEtemcjSXBpORB6iX/SeB6OmHWN/oh6q5kUXC0y/mR4HpQ
bSYHZ392dhg5HJnqQlQNET9q5MVnMQR70WvomVLpvkSiCfneFCIObSWwIb3r8B/x
bSi0TjZe2pt2JfQfjKf/3MF6KAFqsOkwAFzPNsV73UV0rZyFNR6pH8pbNF6xWtwP
ht7gGFszHMBmxOhNoCs3F0h1uu3blaDlFVEfVUa3/bvtN6Ns6+GNU592gP4ZhlAX
/f0PpBXyDt19b6unNVdLhSLUbXRfCFdRQpHFOXz8oxiInbueDr3eUXfzj0HIJVvk
cBoVytjvbYX5H7vB6aeaXxfuEwb02JAfAqmPpQFRtG7ECdqiy51QnJm/aXeIQIlX
ildmkm80Ft8n3FxoUTpArNYg8IgrvIflcEoZUmQPTKFNqd8NU65GDApO3XiMh4NX
AGYbB+hdrsg220GbaOo8kG0gEzbrOQ3PEU5Rs4nMjy+UyRCSCqMYqieU5UnCT+IR
qJj3Vk+B2RCkywXm40q48dmzQ8EfR94reHXNkQvE4qnxscAtfvLOnegYwlEps1ly
1dJPjWxKsk0meQvZ4iNx87LxRmO5+mfMAnprSG+3LgvfbcqILdyweE8ajwhRoGbr
Qvpz8bK7jIfj/tm71KYLU8o73A8Di7+B8CRxEcWIecGdZFSGRPvOI+dX1G60W+kR
y2A5Ek5a+2pzAo1vdUAHgCeIeklvSZifhl7g3vXAK64CwpG9hYeXlKC9lDTIEIwi
Xu3cBLAmtO64qqtJ0suHipZ5Tm4m1KbewXP26fBrNI9Efdarpl+wESjQKJqgTBRt
oEus6Kp/j856FfXdNElSvkHzUuiLO5PcqUOgG7ootOcUJ9wWU+AES9DokqwFBOoX
xt0+FqCx17zUSxNUmLc9LnigwZVSn91AVPrfpAxQ9CKNuDop7uXURIbG2ZzKyf6n
eFmZ5jTudtDlwGUtXbA1OnxV74cyE1jZfkUv9WtEsPVm98WaDHi2EVSO2o809eo6
+SkgN2WunXkR4kabnYkafkUgHEprBsOn20/PoJ0+Ntq4/3rg2657jd4HwhpCoZfc
B3Ccq+XUOMdj6eNn3CeIwp6uIULF75IufNwxDzF996Z7mmRtYWG2Et3KZsez+zDj
SA+I/DK+TxoFKCCxrLU8jH83vABWV8yiOIWzFERozCaVklw3LQTCtQQaSE4vYePF
e9uwVmvtraMJMyBBY1DOcwlszswoBybH0Img9ITzx1DBOc2LaL4CW1eRgehSxXBw
Pwf8BsJOeyfE97cwhsI/oCX71wOd8VciDyFjgdB0WS6yU1oNsmBFXmdohoXK1603
5LEpk5Ia3s/5/6sd5sECB4s+Zb5m78pSws84vWoz740O7+gzAFEn10wqSTDTZC+R
nkLoyvcf/pM5Il/4YsIyWOjlG0ZAgj67ZS9XaTr74mmMI9Txt+j1FJiDdNGiHNXw
DqtyKxymsrN+GNieFtanw1V0oH/CFfR+qn3lz4m8XbfPOb25HrjEiC3omYYCkQi0
pkfq7048h83lv+/1by5qjxk1ZYkHuLK6y5wjlPct0HHyeTY3Gn2FL/IPN0a1oeMS
wq7YqPW22TCI4VFKGXpIxUrK85aj/bkQTNOdW5iCCzU8CJKssZNWNF8zhs03ruAj
XWH+AGU5/99MTBnhFliy4GEjcJcuuP8RjxbBiQTXvqMOucxjDQOLBh4dAP3zfKR0
VHfOgr5dSwVxOGEOgk6YDMigRqoRRR+gSzFI60hv8xlFR8PFrLPQk5cOWXb3qf4N
5p0lH+uaRF6N1DUpRhpdF25f0qPzaVRaz15+0175HO76zkkgpxM95OsTl4AFOj56
ahx2VnEhdbZriKgdcAnPSX7uGVq3ziBopFyl5ieJXKNQEKr4NQIchkTVjZP54f/R
wMVpTnbtHwTXrk6WpJ0K3efUu0G3Rle9iV3H+4ueA3aU9d94MDH+cGIxGDwyqEFo
yXR/QYo6qbe1GuuewbVauJVa0xZ7dHgecxxer6PmcuduWMMRMK547wNtJ9r2IQ2O
YjWAmyioilSyFyJj/BlhW5lxbmvhOZB6/pqSMi4LfRI4nxldaY2GQXTBbXL38K+A
h56ZkzDRaZ8LQ+ksRfe8VjXLVcEZtA3pPzvFuLfkNm9y4CEuSeNt2KTOMdXyeJFm
MWw6wdsFhgh/e5bDcmqR3cE2qieSgtWXhLPRq64+xZF2bZ8hn2tvH7ovOjW1N+wo
/JY39RHlxrlxcui3CbdXi40sI9qjL5pizXE779LPeDUbWnvIu2Qdq5J9+IQx+rkC
zJXQs73Ap/ZvPOhsjJ9wtAbeJV8hPfe5syLCkj8QXTlkHsnQVxs6TvftvwbYjKju
bN+Ukq6X5vAPGfCGwORxAmIqF/jqfLkCyqT1g0SYs5RLpSqU+ktwI26QrlSKuSfz
ni3fEePr1Vm2+gLOM1Pwu2w8ufNNFxZKXL9gTQPrHIQTBR8B148gp8nngrVxDzta
BMV8cUnwsAwJOzsenbDaiifNS8LnBKaTDuyZFKrwqRIL/W2cg56AT00TEjrBZ9WY
KVJS4LNXBYM+OayZ3ERN/9n7b88n1p+5dgryF6Eq7Ax5zYbBlHWHWALJ4RJcbZI+
Q6uI9M+zN/wqxJuISi0fOtUeql5fve/MLrdfyIfppioQ+6gQT4SBf6EIiuq7i4Ug
ZUOL31XI67RFxjqoatj9a5FhOh3jOncYd8u+uGifvBlp9S3dzp4OpHXZu1qifhec
bbX9YyFBQA3aEsFwE88eLmGmIxYyH//gISAut55MLZmfQGCC+7HUhwR2RXlm/AcP
cMntrIG593Oaqpkfw7dm217U+9GRzo/oKbjcSfNXviEqxxFSVMwMT8aUXnXdv2Qz
6w/S77paAepa4+hNURDghf6/ryu0jwtb7rnyH1yI7T0/belL1MmIhXtb11L5sQ2s
Wl66WGlMSAufmioHcxASBDIHy96X2z4vuEvw/cYBxyOiSgnYzlBKmoeYGeGf0yXO
uQR5dOomGdGxMWb8NsWE9TcKru8BhoR9sPHzL2pbp246xFThgSsbw7IEnZxEDa+k
DzfDkBCEF0G1taZIS3nTfVWiMYHUMOQiz6HtenbKfrbi8mk8IPx0Qn6DvUXUae33
PuZ5DDOowBiLyXUnzaHnuNY1lnGsPwf9jRxQ3WtGqC0gdBNhW2x5BYE9goRRgoq4
UtJNnOGbJ9NnxeYqJ1MVN32KyN3N/VOWpEZaXkTDACZWVqy8/EunR1Erf6h4J2CX
aTMcQt3u1WwkkHGWTeZ3kv77EcsRmNdBoshQMulRc6xdpwMbOe9wuoKikmCx2SxZ
wkuplEesDjfl+rgevNsrLXb8i/jUpeLpPqlJ+u9pvpkOro4Cvie+1cSsz8WsknHu
9sWIhXg70SdnQwOJvqDgN0QS88TraUJPS8K3VThTArc51lKmAD54SeLcOAGFExFe
Qo/YTQIUDo/fdrSfNjxZMBbF1su8Bw2rpN8xje4uFupM2S+vsrHXvXYFDJ+DLjVc
NDN7UYLIWSy4lYAyG1ZOA8/d2Iei0HKuxvaJTwaaPNEvKJogrRJSH8WW57+hJQHr
pNRDOFoABSYy3gPL9H+phdq7hVvFuIbkjb5+tvg7u+Xhm6WPJPFQ2UXPbEd4bl3d
lwOV3V+tA350Z21xKwWrqT/FEJM0cfQb8k+36gzrKNe3MXmS3+AXZsdeWgXPgV30
8RhgTZhbQvGtqrfBiYKSJVV6EALT5VjYUYyaF/FDzWoHxLb8O0TSKmg2jJH9n8/l
2rQFTFMwqUF3D5iv0VuNYNSW8ejBdUZmvj+8LoDdjXHx1qEhPo1u4Q9cuNTYfdxQ
Dv5aek4dCcqO6wsqarEYoselNlhYljTa14wf9WHQnEIUhUcBXKhgjjLQL/JezcMP
idmu0uouqtKXXq5XYzcqo/BSRpQjjqcixupDE4Xtc5RwT6AHQQbPQLBqs7nJ3o8X
7vP1epBFvnHD5aWm57d7k8GDMTXG815wARTH1W8il78SBfv+oij5cbqm8RkMJfTD
fVVL44RMHQYgGjHW0JxTSH48RlOCWxIA2/e6zvhXm4xqZVVxVsFoKxpdLByO6b83
eY8M1TakotyUJqhKsk33m+cIMHX3eLJbvrYw/A/IcbhFxMUu6Y1C/P73IgzlSwJz
ljge3bEC1KKB2iH8LRGwlfGhnLgc/U5gmfDqgZB9MlKL8+Z0pEqLdCtmiBjdnim6
VefXHrOISXjMIyA+QZ+k2bBsb76ee/TxgyABBAxld4lcxiGamSk1v/rUeDZW07Sn
v7aP6pZTeKYzkSjf1NQL8bkgXPsTp/WNfy0IY8ZxDH+PtX84S8vbfaq/gBW7xZlr
wV1UpnLtDmtLpjdG49Q6rNYkEdvuCLUPDG/yZeoWtIjJodRdeNXNeGLD2U3JJD0S
EEmiVPLsabAkZB6Adxi+wGAhwqF0jSq5Pq0uBEpMOZ2pJdjn2TW1yfT3oru2R8g2
71kaBhC3X99OTfgraotCXdTwCETk85V0RQgEvsZwVFggdQdr+M2DI/s2zxAg/I18
DyfaRlOVznbAmrhR5snMaVnXgINvPEz00UvyAMPlTn3QOt7k3h/Szvg+eq9TEaju
TMWxE+XosqkpvIJ/B9Ecnnj3CG3G/Us1muryUVYULKf6Zoe1uejdvrbwE+4fC3U/
tNaAihorLYx4zZPxTXKIrovELQy6P/n5UB8uB86XmTdNJICqpt1A5+fdaOj6INZR
NgttwoWL6nF8CoXB50De1z0UZ8BCs9f1yp0gjDIFn9UG5kk3x+WXuuTeun7ZqjKk
Kb3mYsX2goLEt9kDyCtlfHrKVdc0I7GzwMHbBpjECRcbvVZQEmJ6TcqvVKGIMOi4
nBkhMrLBQSS6JTIsmCjEqvpMJmJXbYLdWgVXWtAZLyjt+apSgHijE5Mg000P5rTX
Q0+0VVFfvYd1WRtouXOBM92R30SPyqkR09XMYeBcV4vAgrlndG2/hxoj9cQ5Unyz
mRJwQ2Hjc/cvvGTiF58uXrRvpJ9ppum7UYEoFb75mnlEqz9REu6siKzPyOMnEb4D
4JDatW8O/+JbuoFUQSG+1TlDVjOKbRPd7R6MSdEacT7pT2TLJbwIBQpj3sg+24VB
nMCwoGOGOkjYoUWVYXr7MU2NJU6Akcrjqrt1k0P0rG32g/ONrXCquScVtEmL3YIR
Ab6Y3HxM7WGFxztslzdWI+IoIZh9knknIW9bDzQvo446MYwQDekFXRUNgWxrPyX2
ZHjWh5X3cnZO8ST5svv7lphDno0w1CRataSU+ejtSbDCZH6EhXs0Ew9tzpI/F1T3
iJg0SsbUlbkR9rC0NgSVxnoxqNvoAv8zv1rI+VaHulOOdalMJ6i8yGlTmriZ/BPB
KZ0OZwO9vwp/kgOAtJPNQrwOZkostYNniIqjkBJGm0bh3uCwVN79NqYqTc8KtV75
uUEZUPDmjFiDQhr2FRI+54XI3ierdsJ5wdMqQGnEb41+FKEUR+s2kgnaEb6JxaIi
K4m8zon+D7lIfpvPmmOH95eBtvSZSEl5YPxnmeOAJk32OoDTQ4pXdXbpCxSS6TTr
e0OHfhCfM2Yo7LVX1uRueVODbxSm2HYPEdnQojbv+4wa0RsqitZzafeOdKuokUIA
bgVA1KNQa6OADJRFDBjOB/eJo9jD4yQQK6FDtTWDDY6MlKyfFRQdx+V++Wx2Gj2Q
qi16EKBmKhQWr1o7ocDbX0Z7/PL3poTsXPVDFLMpcLIRndTOEkNwwJaQKwwTAIAv
vmIdwAcd/JEwD6r9SqMZOJW4mTOMAmRjMjB1byJs0/G8xnGIKdqn2CCcfTm07jHP
d0vZyOMHNVGlOWktty92Qb8CiDSzOuhQpyAqHMOLKGVxym1TQCFnFa6w1VgVd4mO
P9CxwDXvZx+Ji6vnvkRRVfuNef0k3IcfTn19+am/r5JMHOXP0meYWCGjt75NtXhx
DLgmIulMQ10+YjblyetY7dKON16CSYGy5TblEPcRLmFv82O2TMyQ+fouwXTxVAHh
W+qPc35duiIcVWT/uS1GUc8biVLXFm2MQJ+To/E//TojuPhj9pw1LWhrVdBXC8qG
GUFRnv8r4ng+g2ts4YDoy5Ty7pMf7OFe4PSRxJxZmKW8RpoIvHQ5o3m+fT8qjMPJ
qgfAzOB39YbsrAAsnAc4iZScxEx9Oz0zbOcGGu4qS0tKh8R4RNrfM+xqZh7OGeZJ
IpJldVN4Qmdenje2yEJc+awnWhlyNEOkZLwdMquWMSUSCAF+MowdBZXJkbFu7TZb
S0lHRWynE86ivdjK9iyzNwyrjSXWRSi0QMkRRDDmjR0ZBU8hF3ad+vYF9kNGXlO8
qE6fs4wKnVBBDTb4Pj/UUQ2KsNvKN9zO/ifnlU0rWEieDTvoH4JPJ1PQlVJ8jLH6
kymLMcL7ZOspVPRzSsN7UjGbjnoUlWsYuzBcanvuK8KAQGdfnw9MyixZwlcB/uDf
nIMRnABAminWlvNvCDoI9ToCJRfWsoZPfP1PNCP/2MGb1bLtjxjUIecZ0muavft6
LAu7ZbIerJQQDlNGWoRREkU3fdQ+YJVYMmme9gHOUsvt6ShqZtWNTvAM5/6Ph+xG
aFAHRJ0iX5ZFEmHrN3J7YB8b5JeHcegL+IwqXQ/a37GZUEXfpT6zFZaK++7yxiPL
P5MndTv31/XIgB+uiZ1gTwQYAutZA+iDE0xhEpJHob3FP0383Vu3w8Q0S6WQojsf
fg0pSgDpXDSgPt6/xBTWgvlCWgjlrW48Zd055ls+X+bI0FG3vx3wa0XT/S+XFJgG
WBBrFizvcg/ofSzlm0oxcEavMJIB+GYIlUn00if7AY4nwajUTOZSYzSUcE7Bok0z
LAJ/5T76U5r96cI8eeNq2RQ0VRB85QO9MwysMb2vvppYd9p9x0xrdUHkLeuaw7QA
3JOOKkYq9CtwbfEcFPGntqczQotc7YyPp9+kqVEouAH0l9GpfcRDbdheoserWfcL
C2WUnykb1xXxzySaILGZIxNXVk74ovj0OmgeyI54QIcUNhqpOHdpKn4ajXCkczx2
WDhmBajY1HHe+WJeR+tXSa0e246m7graavS2EzKxKWjk22GNaZdMcGEY0YsGT/TF
MZ7EahMiBmxLcF1eM6dzbAwvVijp4HQkodhdm+3PjdrCeBGmQXn3UolhLd0LkxfY
v5S++MHeqLXkq8WPyOvGBRgQUfDLoWuTdXRN+PbTplXAsPoo13H7jvB4uOEik039
Xn55gWZJ/AOlFqDXt767f9BV+CokYXMK/L/sdaW89eEokD123tytk1eXY0NGf0Bz
o/lOb7qWjICCNws0WK+DS5nz8Y3tX0Iw9xpg2QpWtkGdyXKVaCiqbnlV5WLldaDI
tvea9yDZWB3EBx5J2ZN07S8M99P64Ekbk/Yt17Va6/KzEMS01OrI139DHBeHJBIB
He0W4IaVloxgRIjKMgane9WCZ4+LkwYTmsETxnCX/FsXfUx//ONI3sdONau5XlSv
qUTkoRDUZQxRYebLoyFFYKDUNu+CpnGT1OVhwBIO6OlVN0U64l+r+13Sa+oDrBMP
I41XMjT+/GUGemrvLaebucPgnz8lnYImAWTkwaq11CimUi4LVYqTZqEAF07NTJTf
V/Go5m8oik/A9sSn8e0yi5u0oP75AFkKyWRCpQLjAz2KFrQeKc1Z9y7c3uBzPOcb
9rIndQ8Mci86Bw9i2I+rDT5Y+fHpUBvzDH/WrnoaeY12DnNgeHlEIXjyJEdEJw9H
Dvi44IAnsOBlJKzzEFqKDV0eW1GRZXMX73zUB++FJVkWDCbNeEKYXMygsxtkwsHZ
8c3tcJ+1rqsclxknlkWJtrwaiv4sb5IvIcefKmjP+7+wqvMpcUDd1iDLDlHx2YiK
O5+4x6FrV9HX+WjDJIyUBoa/zF6z81TijEsVydqABdDsp0GsgbzP9XzA90k3puGY
DX8F8HKvFT5CVYwKDRXHIQVAKD7XeKxKTI1s8tvRepZC8AUV6irQrO4kIeG7NKsJ
p9rke5rgO4qscNIyaSn0qj0Y/24rb+wcEwJjBpWjUjU=
`pragma protect end_protected
