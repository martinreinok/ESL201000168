// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H\3V#;4WDR8(ZM%L@WRSY+;$K^(A+)SL8P^9_J5-("_WD,T.;U1$Q00  
HFW8UXMC&6VA&:U3'O@_3W5I"#_ ]53^NK&[.'0N/$]*(H#&$)K&CQ0  
H<(V8=>.D3SC[QQ"+ZA>>(0I_DB5& 4[QEUA)7\ZP-_!.)!K/Z-D_Y   
HRC<."GNMAB- U,DJ3V\#T@^?8J!1 :"CB?AO&AR/> ]V]<:^!$TJC@  
H*@*$3V<0<:O7G:*[LOK!ED-07)@)COA]T:NM<R"RR"!I(=N);)\V0P  
`pragma protect encoding=(enctype="uuencode",bytes=9280        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@J0GP5(&O4U%"H*CK)])0$95\K,UZ_5_.,K Z;AFI2K@ 
@WQ34PWD.!!7T2F1C4)%"1O<IM$R@DXV=>!RDQ/%ON[T 
@1+_5O[K./Z4+\I,ENK$;H)LH5TY/X#%3.>NUM@)7S^< 
@,-OXYMO'Y6SC@MQ2[I6W(!V5<4317.<&OA:V*OQ6-%T 
@:943H*'9DP SLG?)L[1$%F 5?!I[ HC6_?Z/Y"=96/L 
@:)0MGR<S0I^W?L]US-0%U_2( :R.\ X2#L;&W=ZG9P0 
@L-W7Z(N*I&8^@OVD,W-K;H:JJ7^K?V[Z]XE2=X'KM@8 
@<OR]+>V0H<-,_03]0<Z:NE>.DG>DI=+)G-45(UK 7B8 
@L([<LG\3P'UO(2/Z/^@[OKEK!3%)RX7$=_8@6WSYV_L 
@\QV?]#KHB I2#6$(7-MM4O/1V^=JDUTBI663?T5%:NH 
@6F^I:9[9GFTC*^DIB12F#X:*LBOIX=.(0'O@)+[ZA9$ 
@F/C+U?LS%5)E!^R391*SVX^ BBY9GZ.HI^.P,T]L%"@ 
@_7T]8,]I>_55>)/RX>C#_>9_Y02L?T7SM(*8'HE^]+@ 
@Y25ZC1/]YRA%"9][W:+R-'61;'$.=+ NVH$!"O?[3@T 
@#73A R3]9(0!CA.YEQ>K34 _%B;S_=(;3RP8DQZV!9X 
@(P"]VHZ_A@SJ@L%%<=N?4,I8$BE%@*1Q##O^9F71L6D 
@L_D3G/]C#1.F*$6NVP4S"8#Z353_7J6">.%UAYDFKHD 
@MN&@%49 B/:"\&_'Y;<G.S3&:JUTG,HQ; <"E?4P.SL 
@A8M1#ZR9"0ENLD9>1/X9XV!0H<XE)!797D/1/YBEZ3T 
@6:3"L.+%6CA$;B06V8PT#X#:U&Z-T*N9UPL0MU'?[7P 
@M)K)H.[;N18GAQ,BYGGC&R56!0,%S2]]G5,_%HMUN'L 
@(<6]L];Q3"FN_#6L)N[,^C_/WQRH&!N[-61Z1V%_4EP 
@70R[[:5;B I0KOMOZ.V<V)1<=@2J:@>2&:#FR_F4EY\ 
@2"1]UAXUG>@&1AEM^ZJEZ]#;$Q0<,&?B<-:/?$@_XF$ 
@#IC3I4<B';?2"6O770FSU&M/5>NB(F]U#I%JMY("]_( 
@;@R7)"%:07^J]O<51-;"^T2(R)W R6H31K5=<"JX*!P 
@8%2C"<L:WJH,M@E(A!7.U\=&FG<U,E;@DZR:%8ES_ZP 
@!_'G.YYXUZAO(Y!MT,Y=<@AE#6-:RXY1>HL %*6V#HH 
@3]78\OT4LB1G8R*VP5K4P"F'Q\*AWNT= I$TFUN#= , 
@7<27Q0C8M,5.:4BXSEY@:W#>'TR3;,=+T= #A<KKK<0 
@5<(CC(PKE;1MT3V#5U8-4G!ME?C91G:^!'WF$9_(B,X 
@F/HYH+P2"T0*FT.Z^WD*0>:QEB3@=/_7&=UX<093^?@ 
@*?3'[5_X1[=1955K$E4Q_\"X.Q0PTY&GUOEU;CYO\<@ 
@)P2^I<W _SX8ZF4P(C*S!=6KX+I0)S4P_H'B*(:=5&8 
@^?)!+QB;J5QW(%+-1N-.1U**2.61Q8Y9#W4+M/5>#)L 
@_!::D1,<UA+)[WX[.CSK]KNODWA+F-==>RF/F#=<"IT 
@6,B2)HL\HF#E#&,5>.PEC3H9?T/L\-"?\C9#59B:SX\ 
@$C+@)RE ***-M<2,HD&37$3[G"SNB.IL,%':S5S&X\( 
@K7<G@Z_5"ODDD[Z\CM&[P]2XO''S#09E_=&(</.JR+< 
@X=-3_[*!."3:<<T7\HYL@G?EDN$UK!*@E^6MX>^J?2$ 
@/@<-$4CO-5O%QBC?:0W;+2FZ!7AF@KI&CRL(=.8Z<@8 
@/5W"&CWR^)>#!:? [Y33WUK-+! &7-$"/J]\<>#QO-4 
@M;L_J8J\WT2&_NO/_S[>27'5'GF_>_./%X$#X^-6J2( 
@JK)C.PK24;8>]#( OO4P*L04XSHN%B#%KC'0*S-B3-< 
@A^=VW<55?#MJ5WW456#P] -?RU?K?*&)> S"AO>*A3$ 
@(NOZT8]X<5I$C!L\.];3)4H$7B?QW>06OT9$]'2$7<$ 
@R2JMWATO?&%ZE;%I<,WW]T.R@ (H@O^<,5)39IO?F/( 
@Z/3%K!G8U8/P#<=@JG@!)3(^C!B_#IV>I09Z[T.B Q\ 
@@PV(-Y9/8QH0UK=\A\K4GR:8>A[[>[T %H-O<X 58J4 
@?'CM<3 =LOTJ7.N9R*H;.HH:.;J1\OSZD&6J6<*HU%< 
@=9@=AX*>GK+@H>/A);QIR!,3VKAJW%ZH@0,^$ZW!_3$ 
@9_.P-*L^QO_YERB_D#?[%'1)S-!MQ<L2D?7@2+5OE-\ 
@GAJG(.JW]*"+EKC-A'3#42RT6W\%286K(^?D8N& GG, 
@#NLIK[RZ]E 9!E2N)WRYEWV:QX@6Q]V^1F8C.VKH-(P 
@3Q!7T;Z#*[POB:H\MOY-9,%L0#L88Z)4DSX%3N"C/Q$ 
@)@/YC/$J6]KHY9KV'_]77 \%S^E$ 5R6SWZ5JV1B0^L 
@\W4/[OCY=WKB TO<=[@RT;MT#:?JKVC2H0GG]CO8AM$ 
@%X9)XY?RP\'=C0(DW.H"4C#@$R50@<%R+%B$-:20Y7X 
@"E@7<XHPB L&Z(,D/IH_!+M9[H?FE5&G(B6S).B61R4 
@7^S=J;'_,5WV_^RLD<6V!H83=_L:;*:$O&1K2%\G#>D 
@':;#<BKL$GV@.X>/E;#?X8^;Z3H021PU'>G4Z\C"8IT 
@:?\D585 6VWOUPRU+Y_.6W\N1Y$@%DE$<'Q[[ZZ@3*P 
@/GCBC!LROVC>GSI6.7?_Z^*@+(T(8B@<O>F4CS]ZA;P 
@.\[=)^Z^N_M2)I009#Q++C2^!4C$7NQW_C SZHQ)!E0 
@"Y]95@J7*Z$>6B:+:L8%U&&84>\LE\( UOXMIG[^IM@ 
@4^<KB5:A1/EE6&A:>UL7W?"1W^U5#K]=FG2=?(8:O*0 
@*XZ\['YLDS1@SK75C'C_X&87@ROD+U""O+KD%T5X#\L 
@;0_X=I6'($EE&CN5V?,<.J>^/Q^YJ3%#4V+.+RV$\AD 
@]+XOFXQ-(DEH0A-U?FLOE[F.IM3,2+7DZ/<$AP44IIL 
@QRHS0_UFF\&.+;:?_F"H;H15#+[\/+Q/Y+QKD$,[144 
@\,*C_Q8JJ-+F*E$0.TI=YK!(ELV:"T>1@,;B7J>U24, 
@0SY$J/BW/V'=4.0)?I!)]P2J+E.#T!HY/K^X)G+)2Y$ 
@I]:'4',>CR"@^.JE0YV*!AY)7^YR*D1E'J28%F7I/DX 
@&>6SBOG3=,#8'U^X#M!Y\75WK(KO($%9(FY0[8X/VL, 
@E_5"%-@+=A&>=*P3ZY=T]'?(OX&;F[16.B<R9=GG6:@ 
@6^<6K:&?59+L5@\CI..B[YLVYF%D"LY_UH[:^C:&E(0 
@&B2#]>Y<B#^8(0J0*%>0(N/XQ?<F=C;]X/%("_<^@VX 
@#$2M*Z& 4>1Z;%N9_I:B*&E-?2Y0;D:8Z,M*27TT@?X 
@U:J=:JR\$'O"G>:5:OLVFD&< VLYA3A ZP[!0<HB[8\ 
@TXDV=0@4R>)C*SPX7;20?-<N[O_EV1$\\\<$M/M[GPP 
@X-F]WQ;(.#CV82^94+#!ZU]YC3#%18TVE )FQ!^_YE  
@ FX/RK.L$+DA^I148/^UUZ,M_>\C7;T$510$!5F9>&4 
@!POO% 4LN\+F&0K=WPFH=]JVEJNV%3S(YZY+&ZEE2J4 
@, QXN+8RW"'2Y_&GO9L00!$5$K?/AQ< 6\8;6^:;#_  
@CS^]9R',50_[#U[0-/*F@';(>HY'BUI^3([5,NTS82\ 
@9AX53C-IE<0\/47M2<W%LE;*GFA0_"TSH  &M;88ZCP 
@+&^X(JMG)?0:X/Q-*A<3#S9;1PO@'L4K5J2DQ GD:U\ 
@T=J;KG\1WPS-ZO/(_R_76C:"QF:5_IU-WPK<"U3;@&D 
@53L^-I3\D*=$U 7%(*R2+[.-Y3)S-Y&!!W?[DLX2B&$ 
@ONA16W-]O1>EMO'*PI'BX6TI]V,G0.===9G7)MOE$30 
@Z?:VAX=SE\24C5KSB58Z!%XM-WV2A^I,UXW>#O3<CH< 
@AX,6I5]OK@DT"9XL%\JDM4WPX.TQ2V!X.)ENN5YN!$4 
@'')8HUHZN$-LP 'IH?L#X@7)[')04^46W5M,F'0LD>< 
@WPGK"1ON;U4%E]%L6EMH!+DA"R1!RBIJ,'"0E72R^.< 
@6VL'/;3O#KD\!^:I\5R!U+PG_.2D^TIZP!P)-J%-<Y< 
@$.!@4@M;3"0ZP114]<\5C-AJ R?3Z8<#5K*=4I$#N]P 
@ O\(<&P0&BDF6R3?;K?XOYV&Y4KQV=FIGV=I_;GWI=X 
@+L0\6TCMYC.[;*>7$*&%XM<:^G76+Z4<)SI]LK29*'< 
@\-.M[D$V[M/#HW(];>$M"-Z<X[MW;L^$E5+Q23%QU(( 
@/:H23U16)"D/HTQLDNYI[9DIYC]A'07@$H\&-*L,R=T 
@X=']X6[A^2*FT_3[YU4E:!JSGE4[T0[;=01U6(J[;/P 
@0)*;<^8TG&,@+&>9"2)I!^8?L(JM&:RJAI5RQZJ-[T0 
@QOK$F,M84Y*TD(D7#,:N;UGR+ \2X!E>GA2Y.3G+4FX 
@A<#-S"(%RJ3 '%L5$W9S.*#6=.WG 33PV^R1GEUK04( 
@(UH2H^4P7Q<,D#ML"B1?:M1'1@HTX+JY>O/J7XC#BQ  
@%>OBUP/:Q,WH4BNLD1)1X=*-=;I"HF@@$Q,(W[-+5SL 
@F^47"G<K*,#"S/KQ;2^CH1,V"SH]E$>^O,73/*)+D;0 
@TGMQ(,QN"0R<1&0=&[<7S,BU1H8'(A%_J1\KEU99D7\ 
@.+@/!H4RIN(5,9_H<<^W!8:"9;KC%A@"R$B"TD'@)I  
@Q"1\0+(SZ3PLY)O \E7^7Z6%>02[(2R53A_Y-0A(><< 
@J;#)FE?5GS,4^*DB9@@.%M7ZBVU:@ L@YD ,JL5A,LX 
@:85]IZLO7#(RV-^5+41,/>]I;G"I,P3G:CEKV\,R'A0 
@>7T1NJ\.Q+S $\X$JVYW=@'3UH_+)-NK&Y)L"@ I$H$ 
@P+,#O)D[D)<@G !F9C8&/%SY.K'HC8(IYQ@KE:9 $X@ 
@8$I)5U";<[Z?MX_."Q\=I"[YF4%=;67ALATR_:2["]4 
@1",'$T?(S!VJ=&[[LXA'$+!'C\@'G?9'D [N,9UKNV, 
@M;)^EW6^4W!%^HIA[&BJ:$ 0NR&IQJ-[5"["CE"8IS0 
@Y=(/S&>\B)(XD',36'CC;]G0/V 12IS=,NO$:A.V&<X 
@7Y%_KK"C<L--+56F^;2 _Q>TS L./[BC7L=5V$)-^S@ 
@ P?"R?FP;Y# L9VP24K<<(MI8R-> H/EFLDC>>2IX6( 
@\3D??)9 @5*=7T8()T-JN/:I;%RC1&/K-M\#MXCTSO, 
@:5:%H"\E#:0)$<^PC3EYKG#T2EZ_^[@V:"CG48AD-\X 
@FB3MB11 -\$>BZR(9J.A=*+RM /\R&!*FHH [E]NHR< 
@G=W,EGR-2+0Z))BFGAY);8"3!//Q9_G^H[O@],['B(L 
@.>6<V\02B'@'O%+@TRAP.;FW:"T(MY\*R(%"B\I=!NP 
@%2 R%WV*D]&$D1?3E14=?Q3X@/+<S'E)"\ZICTGW-4@ 
@%T;5J!^-P39\,9'7%Z"6<*E6GXIN^B]'N[M3'MQ-G.0 
@8]35@:W?BB3K 9-[8"Z"/Q)B=C1.=ZY 3@GOZ%)U^#( 
@T&&YR.9CP[$Q2"1EK4X1$#WV3[L MXE&5*\(KJU8^_L 
@>1(@U:.U$'@L%\/BU>XJ0.VE),=U; L6CX.1:+'_PTP 
@-,BB/9NC0TO 1XA,<*Q1^I""K.=_SOQ3,0'="6'U,Z, 
@-Q2C#B=%O>JO/VP;E;W>Q7N-$-QW2\H3^^MO/,CQ'(8 
@N2,JQ'W=F^Z=MIR%0;7P#23>YE]Q-FK\"?941_544TH 
@,8&,N6$X*;8^-0=I^8*8_P72C9UQ?J"J*O*93"N%7LD 
@^3:(F.-^FZ?T[V_!F;%EY3MJY'.%BR -?SG[W+E"^J@ 
@]#$*16!,5D7U\CT#;*Q8T+D132Y9?@]VHP^Q+N>>_1T 
@H>R.AJ7[4W% >/'?P1^QD@=5 <>(Z8-XWA*UY6,^#K( 
@B",$[!E>+IIKB]?A">JESA=M<HD?H^WB+9]2#/X.O]L 
@158#-O3X8B6P%1F*%*,32<V0W8%MRDB$=@3)-#X#Q@L 
@2PMU:P?7;.P(>&/4=N[>V6N(NN30NYJVL^(=R Z2L2@ 
@EXVJ;  " #:4"^#V\7G,QKWEL>/[HKOZN:^&[^5<K*8 
@U;;#D6[+;B$A+%BCV+3_M*87]M>#T.SJOI5[4B#O;N@ 
@K+#JC@1:XL+L3&E\L7A?@ZMFHVX,,Y41NW-&HB;'BQ8 
@5)D9O..SCU(&F0V"P>D$=7Y$.29VNT21/.C8O6QI9B@ 
@6[\/\-9 F9+4I(_4BQ3,> = ZSS!)@$C?'MAD\UF1^< 
@1;6N%H\%[&JE!-5[\3 IBHR2N2ZG>E\S-#)_CX$VI", 
@3%B8A.W<MDU<(<WM/Z]Y1+W!12<XJR[*;R,C(]?D!C4 
@06$;MV%.@H%VG-1D<5\[@133XJG6&;&6_#/O.6A'ND4 
@_+@]^@T4YB#:C%FP6Y,W>XU=RR X#.Z4-%8S! W$C>P 
@]BE/?&:7N2(\19NZ2H$_(D*LK!.U9SJ_X6+W2I(:O4T 
@V'_Q%4DH[UVZ"6/2A&"R<ST DBXF9UR:A#!>A+[WT'4 
@(@-("WQ>1LP7B;IB+26;!P$"IR,Z&]K*E!Y+# C=]+\ 
@!=&V;K0M0&.WACX"D Y><3E)VE:XO[BXKE2:HHVW>OP 
@(V]9)MCB-J_^0\5^<;KCLMHP_@TO(AV'Y =;<=XPG7, 
@4C>E&,R_)(;DW6!&2[X&B2C\BTBDZ"QL<T)*.!FR%CT 
@66I,$ZF86ZW)X#6#98!4S8*?=PK!HL69,4;N@Q#>G+H 
@7S7B91!V<BRY5_6]A>5!80NA,NUYWZID\*-W?D&2V!8 
@%C>I??S?8,LK<FWW60V(4A<U42U63=>&8\;B4'!W4]0 
@26H)IV:0,1/<3#L;SW&RD1"5(?BVXT7=]&]LM'^10=\ 
@L8/5-Y7=2^%6Q"M:)5,!=R&/TT3!.E\S02MGU)<H<<L 
@*.5S,;K"L^R0NER?]H$N0]YQ5'AC:3TBL"+C)@F]OA, 
@^$P>^SY<[W)!#I-^C@,N-E5,_/XF@=]WW0P%67,^$04 
@2/ 49TTG%PZ),Q])(85#B0\/:'5GQ/#NS_0Z:3*9/M0 
@+L?_@@7^^J1CI\KKH)&*(_: DHY#X'JO00?8%=:G$,4 
@X81\90W:++X%PS)BXL9%ZUIA!W-QI/9O6$9*SUX:('@ 
@2KE9*F6\*B76<PM3VZ ;Y[<ZO_]"9OF:I78CH+X\3/T 
@K@[>8Y.@V=#IJ8:(?2_>.(M?*@><*_!YT\L.^:)8E=8 
@+_9Z".%-T)U*!,CZS_<^TA8'T5Z Y9D(&^ M\;5GH]< 
@B,)CEE>6&@6&E/9]&A3@3 &0&NN'^MPRM)<<1G9&LS( 
@+_;QWN-]HVZ1F$_RBH>E*9FT[O&8U:/8F^@L-ODPQGL 
@6)4?\<\L_#/[(,PAU!&44*_#<RJ"_^[.)VDQT*V>N\X 
@O.WV,QC=7_*?K'L=H+Q4*N0>F+3#L3.\-@E^2O^E6I0 
@;+RZ:3THV?0B<L@E&/IWP07P:Q'N'@EP\SJ>3F!QPWP 
@. ?M <YO'#JL% 5E>Y$S&VDE*F4FGU:>OAL&":93Z;\ 
@8!YK%K].KU]NCLBS"L.&]3Q=&"#6XO'SZ,AV4N*W97< 
@1#<QLAM5N>M6U63E$JJ$9Y>OE2\$K;;D5&AIFO2Q5<4 
@O/50I(J?F^OGGU'6S \@LE4([W9FCR7.GPC*ZX5;BW  
@)F=KX1WEU[V77?2LZ,PE N5/>:'2 W+%HV++82R;97  
@QY81A+$E .!(B1J9PDCQF*!D771NL"0CSC4[ *(ODWH 
@4!C%6I(%S61]54U_*"E(7/F^+O80<BWO!? 7>:"/^7D 
@B=[ 7+:GKG>-;6QS/=+$CU(AG/^U?)TBD#:T$+C+2VH 
@RHFKB"P; ,*1Z.#V4,/="XNO]1.="K+?Z-]4MV5Y/4  
@FXR=[F/[QV=_0R*'8V"'J>YW#R/3][L1!G'6@_OM"NL 
@VWW^"F;!"Z!\;CI 6J!*@!: F\!=2.?TDCY[DVR::4( 
@!1I'LJ1!!!M63LH>AWO+O@&JJY13Y"LF"Y+D?)(WGF\ 
@4'X.JT[8  CM#N'=0 W-<]UDH.!R3A,*_J0]'$@T&V0 
@4$69(E"^A)>]EKKEP/@)#;_TV6L[_KKD&+3YW@-TH<L 
@T5>,J]M^ \CM-5S*M,ZD\VTJ9.''[((WIA.B<:YRJ4( 
@:Z]$]1 HX7X"8F:BISHP9Z(W(;_$_Z)/QL&*1ZPSH28 
@,=TP_/?Q[8K630,O#<R)HGC%AF^OCF<I/TTOAYY@9BH 
@*@"S7[T;)_:)Y)S+?><8S%Q:C4L6 VU<AL$TOPZ #_$ 
@L0GE*?<^9.?[?$Z10.>C(TX33; \J\M-#/N-#4)#FQH 
@@XL!F!NY43(86QT.!!FO>2;D>>;FLZ3MOCN@NBL^YKP 
@NR7MD^-9\N,"EZ6$E8QY9%>((#F.L5(Z%/'=?W^VM*\ 
@'A@I1JR\09[X1.*!!O1W3(>Q8$UB(?V$&K5#OFGUW5, 
@A@5Y?G9BG]%T\M #/"T(GN7)@L4<R><?2:*KH-'B)'L 
@[*DFPXK8YWUQ1'?5REHG*AP,ML=*2(L/"9.0\MB4I$< 
@&(M;2BAB@HV/M0/0&Q/<1T80OR<YAEE]\K_N)ER#^>T 
@34B(:DO'# V(O3Q]<IB>56HY80ZI1KO]*Z" 5UAZ]N, 
@E@_2TL3HS3_^_2H\\1.%YE /)[MWYTIE?'AR1>*M.J@ 
@Q;A3K%$"GD]27*6Y_'$#PQ3DAA0\6W>+='CI6 >  I4 
@B=Q7(Y>MS#5*9A6/]C8S<L^?.FUYPC*$1*1NJPFH'<, 
@X$@')0X=S.\E#!Q/YT&T&C^0'CN;%#C52?@0'7E:@A\ 
@?2,T55P7FZDS*9"P&--+%:O>>*P[8;RR]UEUGSJ>1A, 
@"#*?-^50N>EKN38?1A3&,#N)UM#$7JA%YUSC7"R]7D, 
@,WA1)LIF^I?W1!US-*6Q6F_=?Q43:N_51<V&4L $%(, 
@0 ,<)>9/!MD]\S;I"5?)J^TR?_1H/RFNR%,Z>'";7VD 
@A<>-W9#RD59JT$;TX?[!7XO[5"P#+?5<A3^OL.#EG*\ 
@EDBN0_*B(L$C>&?UY9GG1/$8"J0]<V%&^/8UJ<F"]6D 
@W29:4#^;IT=??Z>//0(,"E,*O"[9TQH(])0A"IL$)U4 
@Y,6S$U^=2*C-5X!A)E*12.L!\X>;Y]&CC BCLUS-#D< 
@0BM,\I\A(JQ]0^4''N9N#3B? ;F1D6B8>]=6N< QH*8 
@?8=O/NQCWEHA>UY?J8R>,"@U.^/Z(S'Q#R#:954\?,\ 
@DYKMCKDJ@]7SH1FG^C2PU*'P=!7U\K@IHD<<.'V7D7P 
@!$XB%Q/??$#/N;XH]3R"PQP@U&);R\A1K-PVS.!OG-0 
@.]'15>UNV:-6K6-F<^-W+W3J?^]H. PL4H"097O]C/( 
@8(R44CU)D'@3!@!E&[7Q< V&?OQQ>)IX+I[$LW(\3Z@ 
@&PH@K'1WP,SCM=D?9PE<B_0CO()1\3]NR1>YMH0A0P  
@\^:^NM/6>>$OC3*NP3@8":+(<L_69Z:)[0F_"K5.RRP 
@>T7Z28."S*/;A&GXIT]IWO1+Y+1-4 ;@%#_MC]>0MGX 
@<OH%VEFQ5P=OTQHA'-T>/6-*.'74_C"O$PU9=!+4+T8 
@U3I8\3!\+3JY79AV-\@EH(0-7 J>:K<<Y230V) = L@ 
@3BJQ07E.6IHJO=F)]74*FU W58KTM9UY@J.VV6D3%"@ 
@)^1NZ?I'5R4,+[$K!MF0;* ZSIL:2[P2@%4Z)E9Y':@ 
@?M]SL'4WI<%VYG0PS_V89M.^3$1VLT.5I,U'1N*-@(@ 
@#Z;Y[T\I>4T4&1C$/Z5B@6R%*@M5!A-/\X(I<N\6%S( 
@0<$Z]%P357 6.""CX\5<>W:@&S8])Y*U5&_U*%\)GR4 
@0!5,IN+G%V0)"]E5]9FR63>GV$*JYJ RWGF.6WCEA+L 
@.YH;":-A,,Q:8Z;+%?<'8!%A-3_0D$TDL?2:;*-!618 
@<6W6??@G,66B<<@ 6M]%>&B$IOQMP9N HD$HM/QKBTD 
@@'#6YOPR^6LF6,D/.*#X?[BZKF)8UQ$)61CK:KH7L4H 
@S9,MVB*:R542SA2J=!N-0%F2TVVTG147.L0\J['NL@, 
@=1([XV_N13G%,MPVG O 2>SM\N!3Y2QAH.,6"G_IS90 
@NJK)I_@K!+Q?;$69BV*+E9.Y[&78=F]9P-".@E$0(0T 
@].=\2/;&Z-F#KZB_L++ V>:& %RZ]BVDIH>'C-5E:<, 
@FBWI&>[(_?ZZZ*RTTGXC;@:6B0D]QBYK,6**4%9LJBP 
@N:M,'=&3^B5LEP3ZQ1O,";V$M38;S$GR+*N#_I1XE(X 
@JB>S7:<NH8P::+-0=Q5;D(+K75G5?T]UVSSFLS(MG0P 
@L]/(58,=G<Q!!_56+_/IJL^*OD-B7/F!B >;5 P?H_  
@H'KLF[B>^T:NF+S0'I\D?WK9MDP?-V+=2OA[$U)O4XP 
@ &[2-^5%00IJNJEE K&\B%W*;QB?M6>%X)BG&"'9RHX 
@8W>S'T6Q<E\G#[2\@,NZT#X6? (O+A^5S26:\\^N'L  
@YXC#< Q=UR\#WX'')$&4Z\T#9];ZRNU-.<=<FP4YY@, 
@VO\+53U8C&@]\D6:G$V-$%D!+0:S(Q3NT&D"*R#4PF< 
@6'LOW7 G1?'PQ3C.H2,F80\BI6]!0(EU&J,JL=+K)CP 
@Z)01&?\2<A3-ON'[;_9G*-O\D*CBG_AK;B$,/A_NF;T 
@9P)'7&7CO=/9Y09CP;QLBDA$&.UH4,JTANAY"$YETZX 
@AV.:>^R7J@(_D<Z=5PO]3!T7T?0,!0T70_%LU"R>N#X 
@:T@F&S)RWU_A@T,GJ(;)/4_JK\C>[[O4]EU=BZ4;98H 
@^FJXKHN75YB(A\:'M.5$'Z+-J1 21; PQSO3Q;="A+L 
@^C+&.3DC('":]ZE*-*:5,^VDC-TB; B@:S72%FCG)7D 
@^&$3X?W*20G-]BL=>4%'O,#8B'B7;5" S W<Z*6*PU$ 
@/^G5!/&LPBZ'") WP=;/HCY]EFAP<)HR[.%80P"AZL0 
@I\9O"5'K>&$&MW,4A98*LW*%P>R2??[M4.#5$-/"UXT 
@N^PO5P?4!F6(U+Q C%!C8,0Y!UV3#O>E^&<IAA=+XI\ 
@UX!X_32S%@+(\A$F5<S'E;U@R='HZKUUB9H^HI% T[T 
@!H$\GV''@#]-B\ "#2 W],/G>1XUV-1/N)K5V[4GM3X 
@'9W<QY::>B9H&+%U5U@2X"RCXM8H>"_&NQGH$.V ;XL 
@G#(8P0\@F%E)=F?6AJ@I**2MT'L2@)T)_E2//[@B/T8 
@6;?VFXK?0!)U"EN+*;,&\=/S)Z9&  I9UWAC-QVJL$X 
@TNB+5P4FX;DC"\(JS$!N5D=P:?:9F'(O9(4'Y7Y;5Z  
@@?LZSLK*;4]0ZD]L] WNB0S73+56[98Y*/6C<QJOL@H 
@3W$GU758+\&&N#9O_9D[4QK,/2V(#Z=K7H>M*^!/A/( 
@<C?X2_QAUZX5IK3%7R]_!7%35&SHG@R=!SBA5LZ@K<P 
@B%M#7%T IPX+\4*3E"A$I?<I-_ M2&0N4 CTQO$4U.H 
@0H6CC+ 0<$XH,P4@VAOF\)N8Z7$TPS="1F[>=55( 64 
@0_^K^/ P[&J_ U?,H)/D/4\U$WD)#P 2]&9BQ'%_=[P 
@N+LVQ,?!O\2_2JC6Z:K?+T0N", H0KP1U[65+6Z<%#X 
@^C_BCK,C(B1E6\NL/%!D%UXP0]&-@,Z7:8I1>>S1N#( 
@<%Z_(N^(LO,IZ*,6*$P%L&=O0_4$J:-78@Q=-4)A4$X 
@G=D##7S97_2457S/ )\GNSM_P144U=^ #G3GT1%]^ST 
@D4T@Z136<E3UWC%(RC!2K-\?TPQ?!V7LF.E#'%>U-4T 
@&/IR)5PIIQ\0FE6P4JMF]Q#..?II-.+>@3H'1T=-EK4 
@QHVJ-VY6Q0H#>)JX_M-7*#LI667/48SF3;3S88=8I^8 
@+_Z@V>B]_WBG_IUEK"P 'CW5.Z@@Q-UGWG.^L\X3ARP 
@RCI#(*:.5]="1098U+9O2IH[ MD5P%#D_UF8M32C]\X 
@)-3:>F$[K;LQGE& 5YFK2^"3M"#?@*=NU&>/? VSRUD 
@06R08@G$W8!%N- MT!=)!.?\%6D5WYT;*:O**>P.=,\ 
@./0@H7YRZHUZ;ZS]X@P8:>&GL"\ AF9I+&G6UC\?+<\ 
@4MAP/LRM"'*,K4_P5S^0AS=@0\(<<SUW;-:M+G 7"QD 
@82VVH8+%&2.7\=A7D>]Y4FM?Z00Z47ZSO/:1S-5$O7D 
@I3W8QCV,F2*"^/-=A6F4)BXM""G7T%?RL(8<US/%F=@ 
@NX<5D% K4O<H]DOEJU^U &G;OM'O]V>Z&-1*:L^AJ)$ 
@^C3@KPZ(G?+CS0)&:C25TDR45(U8=XLF/7\>A*AP9-< 
@B5L/<CIRI!V89)IOG;^=^1:S%BJFAH9]E8>[W"$N%Z@ 
@QFX\-MK#S[PB/(+P$\AOL!.#H'0>S_&+VY5!S? /B&T 
@*LRR/%@OR; $2V>G//E)3"M\'SB"GEZ.)O."JD>L&9< 
@)NO$8O2.F A8R/$HR=Z]Q7T-H,7&/XM?9PMQ\H\QN\\ 
@JA40O<_X,_.*=.P/BV=,_86TYA$J@DBX*5%?J&2'*U< 
0!N6AO=A5P<55,<;-\45@9@  
0I.)7IXV:ZK:?HM$#M>38;0  
`pragma protect end_protected
