// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 03:52:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nppHfnRbNXQNe0mBjO48fprv5RjpECuO4zCeM4OpsGc1g0sDRf0hfEIulX35q9ei
HkkL6XL3bPn1NJ7cYp1RDEJuvM/2rDmQcs9QTbK6VPg0Gio5u8xGkZq+PiMjAvb3
NsFF1jFyboX2rl1dq13scO0JB0JvLV1zRrozVJZQwcw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28272)
RGxc7iYOk11GFcIvLTWLnv/Amhj5qJALpUKB30c+VRPIa7WuIRGFkiyGChC/gh7y
KJFYQNmlMpHSWsuoOoTaZ4GO7KTBhsIoX//xdx+8XWP814OxGeDyPgcmu0AiEs/C
CqAtY4hkgpTQIKv1bn2mqg3JznisAswQYLPN0VLl2sS/sCvrnOnHHUn+HxLoyui+
Km7L588dmLZBgd3yRP4uKdylUbZeVzUXLhU6mVHlEARv6jf9hOhiPfRL9Fk/8uaW
WtNiQQB0tvas0CTDoGrPnxA7QMhBSJQmx2zFA2fsShw98SbjBr4MtL/vMV9FDBLe
Bmvj2TOcwbrD5B8agcrVbCMXWstleWM9tzze83aVw6nxkXO+sVBN925dLHjaGK9s
hZUKcyIpWzN1pMA1Ft8HTU0k0nY2u3uhxekyhI+S7eP34BPsKEQVAiltCq/iB5Y5
9iWemDTxh0LVHGdXZ7fTpAb8Y1UCNcUKR8fthJ+x93+baowry05ezWiNOadZfzpB
uBFHhcIUTwD/Ac0i963fwlR6T8pjHMMP9GWZfZwYfezPPQPFUjzc8+TaWoEQRy0m
fWuIkiUz3Hz0bIEGcc+3JfQlEEosBRNo+vi3XZEdFBA6+QvVHzq/M/ALqXc5JeyU
amKHfxsBpJqNOWtoSDRgCARVPRsXXGWAyGBRYvHssQifPwbe9TMbL21v9xIATDvU
U6rLeOHTtUbuDugzw1b8kZEnlN1D02aXJYyDtkaWJIz1TkibN0Dd8RWZSnTAKSck
bpBBcSMi1gmX+/+PGS8/KFkXF7pu8CSqBgChXmQmRRB7ASqznPXLKwkCCllARMXl
gPsQmUgl/I/4FxrOLCad032qE9FMMHxlRqsekuRnsgfOPJ4DiDieGWb/j65k9FSV
hMM4CHZE1UbMhXSBCabFkyc2+tqt83fgss3dY4R3Fg2QJLamw4CR7ssyT7FwCdzT
ArT/1GZ33KsEDkjYjY3nFSBuIprotrMgFwC/LwbfB5jK+iT4LVP5Hel4epjUhwmB
tezRIO2nkp6fNmhhywNtkf/XWqoeTPqfChGE9+8nW+03C8jC+6hhlWRnskTbOQg3
3KY/LsmRzVc79gdDAEoIEdMVkMN8c14PRa7wvtO/FiatH3iwGeRMVK9NYopGorvW
EKZWEagMa+EdklgEET1mFsRc+wU038qOdc5RJfb5dDdG11otocVpw0I/BI+3Qw4B
mlSE4WdJnwBPXZH2Gso6cSU0ixlPMN2tuogl1o221ZpxjnfmYdyaZLoCY0KkVUjd
7LOGHTvT+oavqHyNTo5AY+g6mlS7+IFfhaW7GX1+YvH+yDtTG4GL1Uy1Z+7JgLlX
NFRQ857XNefYPRjeWSOg4VOPr3JSLJDuj2IFHldEnxfmg+IITDN+Gz4jhWJhmfIB
AhXpa+I8uMclZ+hSiqPctO79gx67jz8nhgJNCGhbYmJrHgPESNdHJL16eE+yDt6J
MCqEYh0kD1Wo4JEoOxyrg+HIMt4xrfvkU5jv/skYg9DcllOWfvfrRDU7yV++EF9L
hB/HEJpEBboMQhfTrxWr/vt39b1Uk5kcXzyz3HVaB4lvX7AE+ofZnc196C7Hpk/6
d08LgqJqfWoCx1ZnEuStgbRGILEsIjsWVSp/R2mpOBnAToK7trtXsgO+LBRKEvcl
L6zIN5n34hwnEJxArUQSb/LoxVl9pj7Hx+8Y4l65y7KzfebGF+Det4qUUgIkmB7J
keLIcbsIsvYW3MlgXd4cVJfn95f1cS0ElddpBUHAc7PM8Dn7NOwdUKzSzSVEUgC8
HkT1TcYlD9yA+ixTN9iJhaaDyIBJIJbuoYpa+v7JH2vaZJOz31lU6FM0QjV04tT+
braqq39lZ+MuYOwkoOG7sRd42zrA7//bCwHjBJHDZQ/TesCLTHqOKi7EXgCm6LL7
FKvFDVfVIRkYX0nnH1auotFFCaodkgbQIgqriN6OtXeQeazs4CLkaYL1gvjN/h1s
kb+W1Wxgb3q3vN8oYOqRqWcYD+RzUgoi2PJZvNxikOQRfqjAUc3uqAVoF28BNzwc
lopSJ+nwXpeg6lBuwiLFxLkjKpfurJou9mRmdUGdSYeC9aM7Z5eZb6ujXlCXUopE
VLvbexgiB7zudxQDEQlw5eSS3jV2jTA+Dx1k6go6Jf5b3kzqYD6zjIQuEYhraBvU
2rxQiNV+xHfeEZUsQJQcqFGT39G2iSXsAjAZTReW3X7aXqvp8Sf917Zn6LShRK/k
bTctkzzwdf68NXYMh7E6q562MmF0BeNslmUQ+NJz8TKOppexBpZOMvcLAf4tzFqa
5hiu2CF9AbZQxzVrNpzTBEtN+Z+gRGKRUaMk4IS4CzKsXCJ2vG9n6JJJspTZ8+a/
+PeOk8PEErbCx1cn0NR1JgxbF6z2fObxzf+P8eEpiR6+A4fu7xO8kappM9UlXcew
sq6BpgltYLUmAA92Bd+Ho0jUSmb3ZUDHT7HWD0QiMet4plXZjXr3IcfMXeHnWLqa
sglrsorCOfCb+bOHk7LfYMHToK5sG+isW2Vp5qzLPRSnO/AmO8+fsmfYgZIBBD5D
l1igR9bblaCJuDAX8Jz2zsbULpGgYw62bxUufHoTC9r0n+bH4q4wcZZCJRVxRMr3
OXFrkTojDi3LR/baQ3cGb0YIpfZ5txWpfbt54t9dUulvOqxifp1NBgx5sjxC6Pz0
/gYCO/E8dlx2VXxqll5BkkzY8oVwaQ/Fqt9VFtDz1TG6liKA7wbwTo7/wUBMfOpB
eC/7SdynAR42u/6hSCkPcl7BehYFXWZBWdAwDeCI83/B8qI8OBPdkumBbJ9HOb+i
hswgYNZj70b3YjYkbGmFTa/aBCn8NwdtIF+EH9JsAuMrWp0OemBmiDkQ+9SM3jSm
uNvzNDVEFda9eeQP4lLH3LWFLU+DQhQnc17SmjAtNR77mRJDy0t0Y+yeU3jBtJGD
lvZvMjWOt+rlsAQokrsOzmZgOpsE1/ux4FLbXtjJGB2ZD0SjTlCJlrMjXtOZbKZV
yFkodWdOAZmvDh4YwsNUXJ6IeyydfP4zulkG2vv4b3eHevB4dG4/DJWhdTj6bkJW
xeNz1b8l+Nm0n1U3efskSuKQyypnBri+SvMmNEeX+5K/0+JzrEQvD3IFCUH35Voh
ZZ1+3xYJhOJSOlqME27KlxdLuFLf3gFIigr1z0uPJRSHk3cyxsy52qwVfArdJwhE
le24qc3RLoyJfe65WjJvrmIUexLnV/WkpHhmv0H25cekkoNze4DeV5nUp1NcifNH
EmEBjERZ2yfZPUwDGsl3Oe+J+aaLz25UrlfsVHjkLoR6Pmq/NAPQB60iRdjO73Zn
5JpT74+T8rkgcKZ9pAlFtvxh+n+BJQzvoi4XLwpwZVZF/rptnFy1WdJK4440JIP7
OEDgZuLccInpWlR35yfqDNCUvTUPnO25YCI8PQPSbgZbL7Ai14Q7r/vQNsxdjEZZ
wuSbmSK4E36QMPArZKTB5qvVl4Hb9U0pWoaWVsNT2zfmsLAed+2fe77ViA1aucw5
ALpEn2ytTcjVqApl3GM4UG3XTIKh5m6SYIz8YhSlBiLJV/sb34aXoLVdgBLgx48H
a9T24tyTynr4ydj9fHfi0Vs5eoKDD2GwfvQZ9Lh07S4aPSTiP3rIjrzkpPd7MBjW
FWztjGCg52RwPljbv64epf7zzUeksPRUjwUdNgPPV1E5fEKabE+BCYlFc4uhp4jP
WPQeSc9eUpK/0cHSBRJyN6cDc39DkH01L6nW/GN72Xjij7Fv1cuR+xW0J+QZsZcF
OuOhNZDB8G4K7GJd7hZBMJaXROuepy4zmk1PS1C+MdRdU8rCgQ0cQM1P8jO2RaKW
1GJQz3f8yL+0l6QVGLWMEC6tttEWf1tcLjsuMUy2S2lnO6//n3UD0vKiPOvTPZZM
RCiQ6OkJqhucaUzVuleXXP6JjOQUAmkoErTk07mkrQYiDMQD3TKPpivtq7CThOxB
Dc4iA473yOR1liDAhflaPnOe2CB0I7ihnH/AJ3VWf5WaCmQM5AD09/EySPSLPYiq
7aorzjea4UrsUrBgaWEzQoRNmuTL8yuSL6taxjWHi19J4anwKcovVtRAlug4l7L9
Il1hccMSJylyNBeWA+0+H11RWStD9cGDAjQTk5kVzvQe5L16IkqQR+RrU3NU5WkT
k8w2R5/3PL5r4Mot0Jnl7LtE7sO5HnBMBB3T8M+2X33hB5BpW1pBp3kzm9nXIl0x
GmGTVAzHM2m686cTNn1+m8JBufCOJyNaI3+qzruQoWOwyeswX/Zu3rWGrzHnnEyi
fU7hegwqMIzTeQs1RTAdVxfLOjcnc4ljmdmgocIOCeHUUcTgYQ9e07plZM8rGqmJ
R7y6WOY0XBplrplXEPbtOi7k11WOkxN/VsF+Uu6vitQJEtGV0rluc68Tw40VfWwH
3xaiSFTO0WongBsJ3TDXgRrhJEPnWGh5Kw6D0Z4l9vFGZwmDc1yGh7QRNW1tJ9zH
wmNhm/qXH87SMQHbNu1nzhRqKCkfsxSzm8c9Y8sHkcitkG9n1dioFRvwOb7cS8gq
sKN9T3WWmvulbaW/LeBmbkaN4wt9xKA0Ztl3TzrarLEeSjJ0q3DzSUALkAhc030q
5wsdRKFLtW6YfPvmTdjN8IcPTreZhIEcoUAnyfE1GOndtKnD5i+L6Vwoy2Lpx9kE
txXqupalCAfj2+t1ZuIeFW0w0PlWfsQA15Z3MTDrhUDRapW9hcH/QbRt5DZl94YJ
JEfOf5K0k8oDFxYzTgcI8MCD+/0jQPyfkicLiIvXBg87XjhWAebxVK0DD83xEbaE
cHifGYIuy+Gejc23GhCDhzd+tFJptHshgZSD427K6YgsTn8o3jmEr75Nv5I8sZrd
6Hx4mEz/iyir+qXhkZSy6sTZZzYH2w+jVRJDnyLV3DZ0QJz1V5B8OU22yPviLi1y
uJgvOrwVlhlb58Gqh+dzAVA1u3U1+b+q8H7wQxxJYVHV3YgE1+rxNJfs2+F2Xnsm
jxKCiAX7b0F3SaQ+ph3oANTLMsSQvXTBYZtEUy7nffKtm2QIxOgxh2Hia5zydtQ7
d+9zbHaSmnJGYWvWfwsbmmXhwkidf2zSUbC1sc9GQ9gpcSG4/1v7zJWz9d+JubDe
zFXf7qYoaw3KVpNG/G8ZQJP7V0cIFpPglYakAwxQhm54NxdeLa6QWae/O9LYTe8f
JXHZwnibnjtqRQfBHgEMIjyxgmma3v1DUS0YMM5J7JB+rjWMNdx8sqwB+bnv4hW5
u0l+35snyfqim5mxGHrOIacJcnvWcEKz049j9lLWgCXJR4JwnU8Krmb+u2S9Gvjt
WPBKotNv0yNUMSLivS2McFYPH0SmRyvvs0iQ/uuV6HhLYYtm+eMbhkbJ6XWIUkaT
M5uIEKHFzwRBfevK434Au/1ymj6RtD7CTy9alklRYz0K/bJCP1wl9sUYHSf5z3ff
v59pu30ms7MFaaqsC2OMXD0QLvDaiX5ywfse2+OlTb/EqgaY2hda4js6vlm0YzrB
xGNnpJWZd//pTkF0+6J2793NdATazTmzWRT646iO1ZhjXPr3dsmW/u/TRPkRvryx
cfr6FfjWsuq1wJXxB4WNapj71UHMRFJtFojPFsuY/5IIdLAP/m4I4LmHCOe+LVRE
rfrp0NNB7/fC8fy/iG2anKKImXTxOLGoaXRosQQoI1nH6WsFtEfq24nm3z0ZY0Fs
ZTz81SXm97fwO13ue9TvU0l45+osBvPHr/G3xVwfoxX5ygCdeL0RfvLJDRvXbAU2
bETryAHVi2p8PRPALqh3FVfkQs6nBGbN5+houJYkkzGOjj7edbRpYStI1QbOD7nD
7kugN/jpLzSyTpqa8Jhk/zDoRwuXom7doPZbj77SXHVIp+uLl8JG8NRX2jCxc54T
bhhKsS7FXt1nVgAmgW6R/Z9bFYl3FmGziOYXmidFg5UvJk9XuxICpOtg6fJUWq3C
2UCa3IJu3vSFkL0axynD+Rc1eBN/gGxYs5cwBY8xjK7EcuqWwmlAFk7bDVXo9qtK
gBnYaP94td4XcjauGLVePZx5lR94p83ecLhAUaH/mbQWBXuU4V9bqNlfLue4GlN/
F098ZYxtU39a5oymbThYfrQcCH2uE1iMQoJ59rtnVNjKidPePi/buYT1NTHmzqaa
rJyIawlsKVBrqRoiS963id2vqOY34e7W4jIpbBvQ6nevMJq+tKteeRVW/BJiR2bS
oej6muTHcOFaeF7CONxHGi9YZ6b1Ir2RUqMhWPFW1+sJFSFjyHUGM9DKxLIaIlMq
c4eC1seCpprv4xcYW4/pVXE2Fn23SCfGId3qxrKUKsmF8cE+dS5xtdr7QQnV3+bK
+SpnkI11/NHaFmxTw2Bld740WphughZBqbx1N6CnIACyQgRsPC2Oppn0VDBsS1/v
k7qTtdheR2AZ7xUHKe3x8rRwhfwahNMwITRQi8PRlcruC+xfoz6Uxi7SUk207s+v
PWu8ppxq7ddO/Vkb3KfEPoDiTNajncL12m7CIrnIkfrJ8XT7vno6ZS5beTIrPavH
qUmUcQH0BNX2yj4zj+3nTFHk9+5HMqjPdvYBobOyPOCO2fVfcZKLPrRxkZuCnfVw
RFNq1GqXEE+5BgIwwXHVPRfTRfV8twOjq7yyD+X02BSoX3OJU2usbK3NNZHgr0m1
/q6bLb/Esqn8AmlLw2EP1lfTIVq7y4uRqVdbhqWlmW7wOErdb0T7g8NHHLj4dqly
ydqD6en0sNgAPyNs0C9FnakTWuUQ/hqnffAJsGUsFLA+rS4eVFB36i1nud83/uIm
yRGnau9coGHJiNU0C+KgFYqB21v4WSeiDIVA27KoAcbrlCJUy5E/jo53uk69TwLd
bIdFp0hgF3B00r8w6o4+LrTWotLcsPUwqGxMH7hej+F8u5lfXRNBHAvM/Omy3abs
T53kfoaPRi42eSz2lP+M7x9IQuuIcHA+PDblNy5A1NnGszTW6SK4kl3yINFtw7MV
4eA3Cv7KaTCUGIznDY7eN2/NqNNp27fF9qkfF31TViG2DgaZmk4jgyUJWVuYVHRa
5Yd3Pa7oypZYS82Qn5C5BTiXWUs3i6BM6FVF9Mu/r4oT8xz/s5UmMMV/X/zpZmbN
edK25+YJoaMiBytmRvh8lrz3Dm9z6bPalfdUdmOOYferX1+yP5pSe4D+h8pBiMQx
4CP5emvftdVoJVWCsg1mfwAI4BbRNCmVIs6LZmJaoPiM1ybJfUHGmuyAYfYcjXpt
xovoG13CtatGhil/p/dgHNM+CNUhFxpOJXpjohR86yAgiV7ltnUSdKqnhP0L3ylF
gt9/vX0N8LmANLC/zptESJ98+P+f98GjjbJbVZoH+5UlsE8RnoFq/tKo2pYqrwLD
GxEs2g8Zpw8sIeoSup7tDqQyA0rNf62lGpaqTBsLs4Kq0kvcmfou63TDukkMk7+f
a/HZ8adv4Xca3yRK/d3rma8jZMl240YuZJFvNa2QBv8GXeeoUtwP+bsY0RhFkpws
y2DSoxKUY+F2/hgtv/7/C66WfVaHXTwAqjpHQ2tYU+jLAwTOguJwysPwIftaPJlG
yrRYUjcqB5jF5bTFFcEwmWRvlzbJN/3glHXU7EiIkrwIdf7ogRYMGavL0N3qykg6
HkcSVPueYXt/RgZ6xL9v5W3qv5RagssXqy25MZ5yMSpEMoHUBwqjA18e6hISmLpC
hZulIc4MfdnBEFB9+dDpliBjJFsTGFgnn25LQiKuJu88r2N0xJJzprOCppjy4xto
Na0O646AivoD6LfELpzjpF7DFz0bG2a282r/M9WiFdv8/NUt0JdSyJu7QdTwvgx9
1fnhM5xvpBDj8dsF7CqNkWanMFKEDRYP0jIsIIFdkwdTQWFqE8dnHTm5vGMZK+bf
nxsreoyVBvSHcpIhi/5fXOicYHPWk3TiAdesUtx8i2VZ7E3mxqLKMvpmrGfj9D3q
cuNx3+HxX273/y21NZryg29vJnA3kZi62V//V0fhqcvZIIrsS1Zg7RrHob0GCH7t
Ge70J/S3768wmyHQGNTyNO1OcJD3D/Xb/u9C/8JxCVNB0+8K8njsx1RGwlCie2tr
B1zP/Sd6FVDAjmlA8B9/nniit9wDDvHpPPmjayrGzKN7uLwOP0mlgz6GM57PsexI
9G+NFNXWlGNlfyu+uPU5k/LvIbaL/YET/lAzJHtIOBHev39Pwiyr9lDfS8dpJSX3
806UXO++rFmsSvye5PhsBAahqju38G8o2teN6j64U5L61G+upifaqTg5wyO+DrwH
wVoRnN5LWmWGX9gxBhaAM1sR6BSo6+f1QkxQMw3NQBfkmozF/GJqIhgJMH83jOvz
4v1IUEozYhr0WsUQdl+/cmxYe7nh8a7Zd1e4eSMDYgpYuP6Fu5+KtUVCK+o9FplH
GcN0fEEuBWX6fthRiK29rN3yBFJaj9+g3Nh6K8p6ADeK0fIMmJhcRHf2ekXPWav8
c01ZDfVO4zRzVJmFJO86C4qKeLCiVQYpLEx8Qn3oUoHwuNzArafefFtsOCIAn1ae
ujLwKVZxXYJ3OOHOgJ68yRF6hqklk0ZJbUzBRq5Vxcgb0p+pKJZX+ooSfXYcOYln
X2lqOH4zsn506Qt2EdZkZOHIeS1idWsZGMONTwz/5VuDsF6tSL5iTbv8Ic69FTHd
4VaQH4otGczz/O/wJxvyrHgk/M7K5yr0wjj0TfvQkLPSSE9AHYy6UT3YeSe+MXYl
YFfapKht7FNS7A/nLfGpxAZPqVDuBy7hBj7BqicVYdefD0SGTy5O//Dvz98GnMDX
aRc8FtNCCnoaYOdObu9H1bpGMqgV+IHFZjzyLCzy+ZVn4xPhldHs6Gp40cWRiedF
zBdRINpIAwP5CsObRY1eQR21tTMSbFXTojpnEBc7H7S6Pz1eJE1rOm30+KeXHSrQ
0lEKrrPQJ1ILMIam+hvXdmnYv6TL3VFMyJhgsBT/JFJBz99zsKmgof8uoc+6wpFK
t+sGecNuXpdEF7TdAygPhA2EYR3TcAvIfEUCCHqC9LeOcnzawZ3ZPpX1Y23vBgHZ
hJi6/5o2hyRk0kHRX1PVHEZfR/EhWtNjj5Jux6IKv4Ob5WSaQwatBQf8vRFdBodp
89aiEmNFe523KBiJV8yh7uzLLftqDmn4fTlPhmBxV7VsiGeQ3POL9tQ2kmwSJI3d
yMMqR7MIl5HbmBX0Ozef7duXVd9x3aAx48++tmyFhpiWPjAgE3SfpmYUOAPH7vV0
BMrYRKZ/gmvxCR9H59U2YtPsRqQ1YL2ZL71dustIMkpthqSU9m8SzTRLAOgnRZm8
+pWEN9RblfGayQknLjmi4JUQCTBO0xJLKMeybbCzYuw5m+P/QHSVOvBdQxsSk5M9
/O8PZHDsO2QQxLsChMFoBLUUxvxr/K51Xh6sgAN/rLEjtSpyIkygpHSG/nMV14Eh
MK2k/lVXSF8OCAwcWpNB8MfMh4dLvBr55V8EBx99xZ+L4bvzkO/ZMM+bPk8EKV6N
38jQ4UPPYgKDjKY6oM6FZ5zcSZ8fuVX8/oiAimXs9nP93ye2N51vMbQv5sTkps/y
+x4QL68evCXzyR0JGbgvRs7E1SifRiWPTYGNraG1uKn7a+ibJ2gHkh8fNPM/FgGM
EA1jiQT2nTIBlS+gMBslIrR7oo9JanFkaRU3FyVb/ohC/6YHnlpq6r53+uLVR92r
3CCR6rYE4MYsebLTYhipm76d05yAkplclV4vXVn+b2wMc/TtCFE2+Sj3Zut6uHw4
Itbvd36YowmeSleQpRjfh/jy2mtpwl6HV8jJAsYlMZk3nFzmEKXgBKdWHTJJ8l8w
T7Slu/zWc7y8qhz55+pNFvBynxAXm2laPI3kz9YlWhglIcErDnIArMZByTzUTSj5
v679BbUbMBVoViU/wiaJiw+51xCUWF9zMoQv59ulUFEhnUTrjUFYkcBU9RtzvD2+
D2mMh0R6lUjiyOKk0gmiiDLrilGNwTYouVVAQZRLJp1km9+9fAg6Iv4TU0Rr/sW/
17w588A1d6p2SIQPm1m57kbkDUKpr7IF+hxhhWd/bRk0XQoEjihNsZAb5YRvpJx8
Wf43PDbZekDckjHu6tPfPXCX5pOkpomvxJScwEyql6g6jfIeeMYlCrhntA17aoES
HwM4fyfNUvF3XiP+6L61zD6vMi2YKWYvtwewKn2tofdvkeVQ3s406pUKdS/N8Uef
H0IeVbGnhmNVDUPQu2LvemHwCZI+I/GSolGtm1F2bSvVC2qGiBrlOViLkq/dZCG5
yj8ZOCd1e/7j57sBm0JS4Gt53NxB6Yz1mkJN3799qHG+o5JFGS9Bc3/M9iJxd2Xi
EhaunAicwT9OQIJuKAydeof7kfv8ZH8zduhKYNsW1hBiriHlYZRw8kMt44WBWCLc
mpNEun2OQYejqFeSRFIYrVOXedtIQ7QPlD8VO0KiyHAcbS6FG7wagYHl96Eg5WvS
rQHiLTsesYCaVyAgU1riQAsmnFYkuh9ppscT68/kuQsosdpy5QjrGI2+TM4UdCz0
GxFtCwxYwvkODQrcrAoDltRLAJPsWEZJPIrlarS13h+D8lIbC8m7N5lbiw2H4TP6
9nyhxY6Pa5XiKQcFm1YGeG/aXWJqsuybAWLrnYANAuttXAr7guc5cfuAecB8DY7y
r09TE6HeThVSaazfdwzhb2GuQV7c9d8WkhFUCN7mq6yNIGhB9+GIqrMAPlXUFYxC
rXZWxgI8shOFiGvHHKI73NCg+VTuINJx8hkEaSHdZH3ZneqvabNPqX9ITY+qV/z9
qyXaC2BMDkczCT/0Ilj0bMm0vXAKOWyERdoIlqtOMu9IJMQYG49SQ6H8Mh0TVji1
J+KqD39eX8piSY1COkVU4+/e0vegKpY+qQxxscYfw2qYmUbfaLgytWLROilrOYdz
XqBwCBAI6PEYGS9PikyO5tO1LM2HHQb+Y54b85+ypnT9jExoL72jX8mnuYEUVBBt
5gg//ppjAbWzvorYXSCwGuioQgMr40G+1l0cMQFKQ96ZqENUL2MlbI5nyikvhSrx
GYeMWu6YFvNazTY/mF7EuRsRig919XaJYd9J4uKoROIO1ApC0BILTxkrZyB39KqJ
qz+fZspgxl+Y41xzu/w22o5lT/hnq/U/juAEjBpdKI1iGPWG9Ef+E6doboJx7Q0n
59DakrEiNqjF9Bb0wHBPFJ6lyW1rL1ynpFpZtQha1ZGtGba09evznb2bWwmmLJUG
3+oW7W5Sf8zPFN4k9uOLlMaLveV/WzbjyA1VaPxkL6TS8Fl98xVNL5FWoKiJT6jb
ASEdPLuT/BlZhMuLmUBaA9X69MsltYfL7Ur/JduuBtRYjcpwfFuhGNMToeljpZny
5fzM1HN5aA/isLLed8FXl2WBpaUeP/DKOaLqrqbFb61W7P/5nDkCNv9pxfqHMYFr
SI59RTsJ8+u5DTMgzNtA58/WVhFYB0yYenuD8urLPB9IZlgmtJBYtcNmqZLspaCJ
HyD9sbvpY5s2eOmdiUXl2MV5sPktWTA9l59ILQnIkevvGPwOBW48AvNFrzyUMFYJ
nio6xgqAO+8NDAnh3UOICt3c+UGf+Bz/Gw0mN78/G/QPRZhr7UmWnMbryIq2z82V
hNYnivV5zgPhE0EDDQX0jWrTo32PPut3KNb2i/UkQYWDfqtZB5cUMmjPvyff4tLg
pgugbzSMsTZuYxwlw1w46NsgwO6u2HVKWWdSZRGcxbIK5npl3rK87b/6CZzcOG3g
Rd0e4G0AMbRZ7ciy9q60AtWxhOqitadDCZ7N4nxh5G9yOEWhvCo+yB3nVkLQO7Ag
LBSk/t+LhIUKREs3NYOVHPMVI7DI3Qv3VYb+ja+UmCBrCQ40Jl1kHPt5B2qwGl6G
oKSiyxfbXaUIbqdIOFg63LNEUa+QRo86ewSPH49uc2dfoR5unGLROHwTPyaVj2oH
iphxs80uRjJDpFvfd/hyeETZPaAa4meLMBYt4y6I9mX1Wm5bYjmsCQ10lUCNX2rr
PeGsWzvRGUJ5OoXwVw9mNNgtSfwjoIBy3W9KgcTijkI7q/Bv3k/xNC8UswhzIYr0
si2o3TIJslcq52yoES0nDsia7HXmJeAa/+FT39Eh4c0gwS74qD5Mk94sNbF632GW
Dkm600/bdofHwYGz63Z+fScW6oJW+jyD+veocFVYv4d891f45RmNl+CLURhEczaE
4T/iv2AmY8Gt0sccpLZYCNxAReyu+HjK6pnjpPCHcgOxt4u3J5ncJKs1UepEQ8rV
LZe8niosE56AzbZ+XB4N8OSI101KRlIgzwOwG4yRIN2eHlEu30k6492VLMFrw2ca
FqkrI+KY5NVDMFzZaZXPoPJMKV6XGu4YS37GNA2YZe4UkA7TrxXfldMI2UxlB5Lg
3kwpLRtpFDgUpGOtO4VhQOPrqDdHzvpZ0thwGKngWzxphGnDfWRZkjy2Ch5PWVav
14CB5MR8OhZsAOEgYT1cHtmQ8avl0ftNBS0+NndM/nUTw0+cTqnONJmVksce+DgC
XH+ZcVpiz+pGasmTOIxBTEpZO8kg3RMNnZfBRAiqaz42wi4eSe+CU7bAO0BIYiHT
vVCg8g/YSh9vAKCrK04K2QuMiEdf6s/hCcBBr1p0YMJlDi5ROvZwLcf+y0UEdBFE
r6rpOy6PAwIt0xMfskYPFjNTrKXOvXgx8unRlVBqI87prWXtv0A+1zW6jaobm1P8
Tjm+3VIpMy7pwwzMwoIrEZl3Yigp9M12BjBC8dG176s4VzIMSvSEdgBVAKpBWU7r
0RHsfBXJyDugfuiBpB9XcJ+skZUObtEBS1wzQ5B8EDvCF75eiiWHzpRZyX4ryZhP
tDccmdhmIwO5YWEakeMq7KrDYKYnhifUqPQ0LT6EnHTzARJsCGwVBuOif+S4RmVU
lW9dJg5waDcHTTc1aFrK7UDd+j067CfCSj63P9VuuotxigWi6zWqY7ViCjwG0p/P
CcRlRpxjGGHV7LBptboZFC20A7FPIyGO+BrTyBwuLdNoHwk7kvE5tJwVbJCjtPpH
6o+RWm3XnzqJagqTQY7uV89lTCQmbLUQlXFbAHODis3/VmsEoEdicgCJtS1gAPHH
S74j2lBYuCOtbGjm51+XCWxbtguJgijbOXTxBtBqDHz40tKU60rjzR7Mn+YbluMu
hHTtSlkXmI696lp/xsQXdJ6jPhe69CxuW1bzwnDxUcfL6DfiGXxebTdHXSzW9ibQ
MEgt5S5Xn8fFSQ40QtjtAT9F26fioV3LLwH3Ylnr6y5q2b2bR0tL4P4fAsNmFdbp
DaD+q1bfcb9gsYEayGaoH+tAqMczqiHpwqZ1RmgAEXxt0lRt2CfCq3uQjdtjUZaz
jGzCH1C7doFQhrkP2tX60stwnlaKJK6c+fCeJ+kFyNJ8vxudUVQn+rXizGbaeYhg
gXyStlju+BWI7nsKHL1QGNeqwI6O7fv0aOMZCD5F8tpfRgyH+nWFavTPSzXXZ5qo
PlbBslIIMjb//r7oo+HnC1zHZJ+U4C8v8P7O7OUz5Wt4YEL3/9HrRnLlkEWu1vrE
DBmD1U4uKQeF3ucliLtRUqP4STUUOlwuoE2yqJ/aVNUb1JB5EZ006XG2GWoQ+YUA
Mac+hNSLXjrUpOJIgDR3P67DvuHuou67cNHkXnimycZ0AdSaYChWz6nP14aKlriG
S2k7Hr3P0SMjSqD633Iq1cXDHYQLYqbnhny0nL1SA4akJTuwep3DqPplYbQUjPEr
QvOSeti4pZFj+eEc5XQmpl5kflLUOtDY4a2ZBv960TL/LE94oxyz6n07oT6IGI6r
/HtWfOU4Y4rMAWSwLXhk9X/TXEUc4JseaI8cT3wOnBQhqhrvPBkVhtUNTr/EfL+i
ezDLvDE080seeX+Ljbj0w/ftRnrWmwnRAQYK7d/a2qmydKLdotb1tSfzeRijmLI4
xmeLFWfvPMwuXyQLHcz8Lxq0Lz43EIK8nq83NhKhd6FAHJTlep1bEhkpeeRYg/So
1riTE504gphM7t37PEg19fO4viCd6WnCivUvxRprmHeO/OQCA/w3BDm8TJaNHEUY
Vp3q+NdHR0MhddkagqdV1fltUB38tII75NDGSj8sRVX/nutiFFNTSZOmIyDyaZgi
WSqnS2VV9RbvqZ6zCuqLqKRkVKLPfqlChgn/RkOgik0Y8vE/cSiirX5PYY7zCEzu
5Gb7zQklIC+QSAdmpukpxZPeEYTjFxLKucd78NPYn+ZJ7MmOU1VNUgYswNGzeci6
c317xjhDemDSJ5Pqmr1gO/pfhVzfRZUoRRWKpgLDzuL4D0DZSfXqiIW2Y70JNpdL
8Vprt2cAXOllSvQ3wb/RiNWu8rEoBYGeuJ8/+aALEF40/kb8esLJS92fE+fXTkzn
4m6Rggk3nsy+2mveI1f5bsUEmy4glXh1ig1vOdlPvOPmxDFPNhJRWchLVl1oRjK9
tJX9Whr2iOu5uGgnFnmPEm2XN2PcA3X74kW0GIJQd3/KfpBcA7huZRlVDJExUCZG
PHhcSn8FkuLkIEK51178JREnl3ENo+fs9u7I0wtFtwBqhIwEhh/fPPd6zcWZE9UQ
C5EgwKHKHOuBYLK1wJT8CMy6ctg9T+8pCa7oFbfEAfm/xsYAx3VSm9LEyK0d6DSH
xRIxGcPEzGRCbQruhxrc02x+42QAVsl1WeivsWkxbidRfa7KbUKXtM9qXQ0PM4Wf
uQ7sO2+oQ5XjWOOz41pS316cHNJD+nPpamMTYgRq2RSD3p4oAp/pTYMR7oS4/fGY
anCzoYS+1LA019BLOvbuZPrPwichOepplM63PldnsrfOnZ9RzO2gH6YkZaqTpR8e
/MQVkvHmJc/kxtLLlL2t/CYbs5AK1LBWoovqho/Zz7B7GfYwbGUiK28T9zLTTkr4
iBIX8nzPKDRw3rnXJgfiRwDHPepAxDlY8dcBqmURSY+M0J0Ipj5DmtsUyicW58sX
ybCiGJhOHDPz8rfxIV6VUyQ2NWr0cbWFADJZ4SoP8RwBpW7imgwFtNTzAr/hKELr
DWxCGo51bxoArSVltJlNCIdpYRwoqnC2S5qVVh0md/5pOei0azGl/0ng2sSb5sWC
4MYF4uiESCNNp+Ua0TFcJUn3LUJYVeAXVY8FJr8Tiv27YBOHDwX/LM9iDL+XFA+J
CH7jQFAK/5K9AkpEKWnM8mKrsOBoZG0+7RU2mhyb025ritGF6AO31v7JOGPcoNJ2
Mbdla93j+gY5A0NFubezZY36Kvp89Ms2SGMNnJo5sC9BTBoUj8CVhN0Vq/xApd7l
G7oV8dxDyhDN2bdzfWwzU8Mv1W3k2aANbQ/qJmsYdLv5BOPTcgFfGq3v/xbh89/8
vvS7ixMkGn7P4Bt0vo18+4aaQyKLnlMjMwc2UszLedo63mxgUlTiHw0i3A3THwis
LR8L1Og79MSvD62i2qFn4jehydFt8bzK71RO1pVge8EqUDCKRqVN2cZqhJ4LMMPs
JTX4vK6CVa4AzwdRdsIrM3QKpeJF9n9QB7T5xMvIwXDNaV/imCcq6Tp9W3VuFA2L
QUkftQGqQ0EZ/h2SlPBkunFl6YM2kFzIAVOOmTambM6dnWHYFkLnadvuGi8Ss/72
yUtlEbdS5MH+TbLgLZAWxXolJyfinBmhd8VuEbCVv3FfcOidnhPT2WGy+Y20OoX6
UM/xST/L+iRZwJVPotJ0+bfRShUDbC1ncSgDzZ6h3kwxdddCiV7SdCnbC5AA9+EN
FatcuP7xkVqyf7AbWz0s6xpKwaPFmPM+MRMxE4wN1SafazZK/DLN808J3upE7jF+
LoKdcYwFexju1qHuEFtdKXAVnQJiUjw/QSzrS2Y5TJ5BOHgrlepB0Bwpa+mWwBRr
O4vSIBPWRTi1mUJPhY7e3dGfQGMW0u74Un7YA0HLbAfxdezhEou4Xnuj2v9kl90G
7KvvfdKljLWUVdfSzEoYo5c4kb3JWdoZ5TPe/4VPQMELaOWLxVcP6rzTOL0ldhOJ
2XrrlwA1XLRUYT4ghWxHM7B27NQaLuL7XDHNIpG0BG4L8WyKB8Zxx/xVjaGCpL/e
UV5PfJwD37iEBZgbUWnnS38aH4X/dSigMJP+BYtgqsnKMxNYXMCZ/Stss7Dtkm/q
XYBZbjqGycoKvCtyQBI9fmvaOL5zrpXp1jz+BNtDFYdW4bjnq74UjR8Sii47cxuf
aiRLSbKaId2HHjXCycy5DUzNfLqXlvsqtF+mlUUBXAJpMNVKaictONiw8gS2ZRhR
kFmuYmA6dg2HEbaUV4MS121axWPUMCI7UbDFs9NVyrCrpsKfhEjQEWOh9vi6oZSX
n4pqERxlOhzVaXVsdxZK4oQox6RrooqdZqX/Zpmn4BOTae7+kfv9Ldh5K+eg89Ei
DscLUy/opA4qoSwCCG0mVnihfxsqYpv6Zz5TmJJpuj7DLjAo4ZWzmnChmuwr874c
/XYPcA88RqRUnXon6zwkLKZ7UlspwItlmI6mg3Q3FucMUuYE2WplIOszl+M4MD2F
QhBdEAY+EJVWm0gkpBivGgXh9o3stk8e3zp6QBtHzVIq3KsyedboQOAU0tMfPima
rsh456nhjKz43DB1Sp86O+F1PPHamh2Lm39T1rnUZhu4glnWPX/iqzsVCOR3b7Rn
GuY6sVe1QtREfh691ouhBalVeZKDJ94cHcyUuI+aVljQQcmLIIokNMlmiZcSNKkB
rmOesQR/YARbV36Z77+6k7/Y6ptFzPv009kB8dQq+QDSUZ0P6vuhdxYoho424w+G
X2DQPYSR5pr9JLqK0FonXh/itMyFn8E15ll2KUc89daJ8VeNoUSC+rwzpYGZ2tXg
w+LftcUfzdsbac6gKk1/kD1R1hIePUTlk6LxnLfZV/wzGv2s/QQZogOhc3IOreux
K1TsAQxTqqhmDC4pvw9Vfj2PsvpBYkHOe/fQkAMZkIvEi5ZDiNlXu75Vru2EMUq+
ZvOJY3sSadUioqDd7S/OJM9gqQF4CIHWOljzW2NNOMLHG+LsbVknzo2gttm7cqFB
KG8unOfO9ph8zkChNDz2l/6voEUcSnQXOIZjLqy2hXqwFfZUDft3RPpT5fUCIoLo
3p0L54z0GcflOMia3QBdghj9V/IsAK13dqJBHxbHRTeh5hhELE3IDX4phm9QxAjh
HUx/EYtqskh5Zld24nwcWW6AuunUCFeQ9f3fry3xYpRliUusDiSXIYy24gaB615W
oC/V4QBBmz1NjGOV1Y9ulVSkpqN/al/OI92SSu/SB6HKrkcRhtFmCY/HKrMg0Gbw
1hGcwA98rx7CIApV7ayR6dHEShDMv4cX1yU1nKQNSIFb/to3d4xdhsyDz0Ocs6yI
H1x5AeZ7hBYIQ6AlzV6Cn5/gxE2iAGgviYCM6J40h7sND5K0PhSjIByPdHz4vd2Z
XTbl3CtWKHazvU3YpCJ/2SEA0vqIZx2IeVsqbjnKdxFQpGq/SrcvSTesXnAmkpjA
p9pyPfqoqZvoSTEwaPLkivzFLzmBUJbuX6dyAALx/eJ/PKyDGHr9tgZkz0nZNFfy
6kw6EfRIgwZASjB/6zmddatipKoWRoNmZ8lw4S89SkdSgUZ8L/Vdu/JT1YUQjRGF
EPhhLYKo9urphTyBphFzvxMawl6BB15IW1/ki7y5DBGDKm0COpswuMxEgL7THEDS
WEiZ7TVmkCKBwZj20pycorhHRiOeRHS0iHDshM1E+9y6qPHWM42l9ruXR4XhCM/u
xAU/81g0rRILAShcWmPZ5YF2Z/Ck4dM6uNhD8SX54dxO5i3fM7r1xDiptfp4B2ei
jlXdH+ZbaqXXO1jhkp3f5Jzv8HgmrxU0ceaK/JDpgOPZgj/7UBxG7r5A2k+27JJ4
t3P2KfQutvd0chk/Kc/0LGVj0X0rCpbEtHu4PaiDZXjYDz/11SiUjWNIGoTcSeq2
NoKy+4JRa66Vw1dE/0IPCtZe6Kt46aTht7nPzhyqcP/M0/ySA57bELvShMlce1Fo
4mjIjgpSWEyRP+IPMZlJdtyNGcq51WLX3YSc8VUrqSiT3YPks95UwsZZqpiV60rz
9kquLHDUchdDxfN2Vs0ZI0DD81qWuEFAkcEMbkQWrj57nKJUSuUXFqtJfXqKSzDJ
3zOpcHWEXmOsmmwW9N1TZaULDC9vA0aPquPvLftNiUDUEzVMu4MIj2nGTp1hdrxX
VYrz2ueOfJmjyhfCwt43jdY6CzVEAqTBzYMC1YqqMnKnMH3RF8aes3fHsos0tPbn
8pLDlSibvYZGTeNcrgYLxKU09ErgvrY6fRLl2FxiCtmR7h1P7V/GlsXvF2hut9ZO
ms655ukpHQ1yt+HHd1CfAq6xUCXiI4HULOIhuY0/S9rw/28lQ5Ys1vOdVXKjJLcG
PNsEQhpnAvuExi5TISaYmB2MSDG14SPAik0D251od/2z96TC26DuIO2m/U4Cx17m
qWEV5RLaxariBP2Dr6VwwdnJhvHmKsYHoxdh9NIBMkxiM+6scgCvp6pup6msd4MG
YWYOnbPdp9UMnL9kLn+Feb5fM0Zd7nwQKKxy4hVbYSWCp3WUUDfURJh5SihLpAi7
R+cGkdmEOT2jPfFpzUNx1VI0MtykYSbeBs8UucKrcI3linSvwt7cX1VKZ8sOvjbC
kR2yLa+Ntbogv2J9HQRr6BD4LskAVYwugd81jOL2rkTF0KMzK7cOKUEHkfT/da+t
YK7KWbMiDXHZJzPEjboKirs2wm6M9MeXP0opzuLuOcHonmniIdKiQ/0HPlNLPDZA
r3oexCc/IREsze7zWBuncGWx6v7/piM2HyZqEFNZrJg+iszNvbIQ2Ybk9C/5hleU
fMlTuUHwhR53ijkx8VQ/iIu5RLs/9ldsQq3XpKgHdvjS/Bxp0hY+LfN88clXNEgq
PKREYsRvG0uFapWR33yvsHt2bbZyMJZKZ1lzmQfsISfYjf5cdBJr8SCxpHfqZ+oq
gRW6N0pMxkOEims6YHu9omqnbtgIQyPQC0xAI8nMTx/Nw19torbDHlZAapmmyHWS
rpq2mIR+glizG5yw8ZzeyThkEFUGRpCYV85mbSSFQlJnBOoWP5U5cLLEnUbiaBig
L/0L9ekXPm5QG/NaUjysTaTEEMjBeWn15Giq6+hKpEEkiDdaLzddOvv0UyFP2WxC
KbJ4xg8IJRNhHd2hkMfvhPwzM7bPxHMb526+89cCHv6ItRmj7U5INeKYwdTRaiS1
V8TVWOtiS5wT2zj6tKQrNtNXlV9yTDLUmLFabofG+dutz9MeWK03O4RWbIWoq5ws
EHCYjC+OguKmK0SlMQKiWQqocBEjBY65u+0hVjbAH7Uk1Vdp0nE6yTGG+p9ghr33
Zw8MiyFApD7K/CIBpxBvTU72vQrNe5F82fBBAymT3kQhRjOeDcfSwJ+sS/Axhn+f
P73GtOO9/Wk5o0dqzrn1XroQABwlLxtbIU1iAYIl9y5CkfAHPHtsJwqM8kQU0/ml
pfk/Cf1ij5rPvFKlPbg+R+xFBNtvmPWImSc9mQYpX8rhlphkIA6E3FO74gcIbMn6
FcJVje4QPgXgXtNJvv7/jV/VgAQQupwjvxf/RFdRZSl7LA8VAH1pD68nwuKYV+KE
BpfSuA4dx9qOo82y3IrJO+lAbKmoGhHD96TnSI7vu/VT9D1mSryXYUwWNp+71aLr
kPZfldSZ+JXuAyVsKIlvHtNyGIg/CHXCO89o1IILdlTZEOpp2NzqChyGy5vmGij5
MHWckETkSLjCMF3g0uQVWzkZWi1f2rFjtlHk4l1lDDz9spIbBIDIHJqSKsVK21mv
C5/jZF/vY+LSxHbi8aNYINt+psLgVm5Qa1YANQBWKQqHPdCAlUgakMQuNA5gDlyY
7L6Seu9E7PGqUUftvg24LBi67tcPuNkEx7Tafbi4yWqv2El3ZynKbbGFFCyi+kQ8
pfuIpkrxqBMpmPN008Qe39/pOWsoyJyekptk+WYgnLLwOn0WbjbH92FgrLCSMB3w
FSmBLfrwHTbEcPC7+iIu/zYVuumMgqL/FaGHdFKIYBB+2lTdbfnAha5Cx/vNyOIS
/AkllXPXzkltf6CflBrUUONytCA0oMsLK3CyKpwGknFlXScjKx1cg8Ccewl+iyGi
0r3pL5AR4Pwcy+nz4L2WO5FAEW0oRwLTKC4WTx1zv1221ihH/pE9dGJyh9FUYN/E
R4IiZF+hZSCC+THfqsolYL8mu34Ba9fHoS1j5Bu2odkKo9yOIDI8nMqwps8DcstP
U+RfRfjpSMIg7YYBf/k9xQ1pul7Ra+5mW3w/NRx5b3hIyrmOd1gg9aVgGdZatWHo
ZeRnTK2oyuoa4TKVlXBEhFhs9/XpK5bWLCdKUkVP9F+od046R39iPmnbfyUWP0Mr
kHdBGwR++LOrM971NE5BW066wHITfCmICrQHR/WpM6JvxzHfLP0qKCbgvi8Sofb8
OoZk5sye56tenFX52IXWLwqQ++2pjwp+96/tIPPCm9I7xCCdr3nhqDKF8NlGSy+x
4grFBSUiwKyFSPJZGSoKiEvaBHoY3OjgpvOvOj35t0KNjbYVrWK0Ju01GPsEp0Cq
udRBadTLrTKvjuTvBIUf9VnEEXnUorLcmmw1NNndo9+qFUmtLQiOo/s70wgVymK2
XiPsp39ZnLWMDVV25713ZFFv+VGbRPWfX/RihWF1T9w6Hb7Z+w+xnFARXZRkpO4S
N6YHJHKo9qhlAjj+XnbogDikVi9OQzdgtHhsHk8mYlQA/MrpK9njOXRMTc8JnvaA
u1e27L6fk3StD+OcKPdhLsE4t39Ve3B4s9WFmtEcRJBPn0S5vEMJH9rsRFDS1rUD
I7Lg3+AXJxLEolD9LhP6IBmWTyMIMHqd7Lym/wVksvdV8MuBykaQWlqsW72dYXOq
sbqJfRG1W4zqp6H9bZm5hbWM3IwA3juN945mB3ssXFLTMrkyvH87e+WWPddn7M3q
CvVEifR87I6hS9L9t8vr9FqIgLrSsP7HwijTWf87xQrgj7YzA1ImMgLLGhIm8+rT
sfDpguY6RHfUyNaHeiO1S2seXA+tvMSfv7W8pzBFZPN1qCfPgDSpF0sCONhAtt9I
iIkOq29835nCOsIi0j7NkKoDOQ1WJ8BlPDAij72mblSG1dnzC5+K9fNxzwjgPtDn
2pZWxKf20bmnRpcIlTToUI0x1E7huYS77Svgc4pDlEIG4KQxggXSznqOn+sRtFYc
OpyxRHLmqHDJIJlST5sKgnJJqPA0awBZ4+fWYcWI+7bgTDrNWwr3k6TrEB1rIsyk
p6N+4jva6tPFDSqbkMP5Y43FbbPINXAaCijVoAjlI5rHEWQ25Voukth3GdoTNj2M
cbTrtjaMRGay6RPihBbLOmVLWf72BBuODswz4VCdQj2v9JmYmbPoOhrlJOALb3KP
/kiK3bM2H4xyH/x0Q6rilhWVtRGXVp3/+3C8QrHeKL1w9SHv9++/7RFkwJh9uKOG
77wdx2r6z5GNE9OX7kWpNXVRBWQWY0XL5C+Roqc2xKq2gv5IZl63xnUf6CKyp8Ye
pPm1BnbWsVKoqDprtZGxI9c/TQZGYRyQHjGmcbJOmAwAGT9yQdAUb8dWOrBE9FZ4
4UHbstHO35GIf9bXDy47zjyAmjYghik0j0k0pwXX35Dkmlk4fMg1ZFcg2VEcmNJB
7E6d3PdnoBUVzW/hA+lJmJfazy2Bhajpa8NcnBa1kPT2AUC+8dBLzepHd1S/7pRy
zmjipmXrsJOHSK1bDymnI3HygMYJSYhcYv66kuk9MyZXzyQZeq/8sLJ0LYtPxShv
UCdr5edNrKyokWMmsWCFIwDrs0NztT9VFMGdDbI3PPvnO9DqrUVGDWfGK1ldVS5y
XSdXVE+Lft3X8nRT0y0Ji4Z0n5tzkeDOJEr6IL/+VxaYSUqLvXZVCD8NKz4sR8xU
54U+i/i7HiARs3kx705579plJe75zFHmEiAOoYRsrd/KRzNMORy4SZM0EUxFnnKr
DteJEUgVRYpZcblHUt19xodCKvM3Qy7m7Fopb7u6DEPKrmDDb3hb3/+pMq9mSOak
kKDsX2VRBlsAEW+qE5vCo725Qujt2Bevi+a0uXOTkaANA69WL6Wur2slx70yotty
N4y/Nzlqg4W+lCgkS7RVlinc/gw4zZFEgA1RtmtmVWJ9vuY5bS64eEHIadurVaR7
fa+4QtMT7rKGKTyBAA7UKazUIM1tPPthHVjjgudBMwilAnXAtpKXsb2pU+OPqJaj
M6RsBg8iNth8Nr6xx7UDKJAnWKgPptV3cySB5LRBiGrLaBz+A8kHwTKZejdkx5rx
TAtCsxPAuQ9qlrT4dOewTPQwzD/lie9Ym93PivpC+E1Hcp+NGJw+aEGvK+kjpuw+
q9tDsBupCCscENZhBO5jQ6UDt/8cQVuuzOEmFEke2LaCX9XvoG4wkDGjgsXd1Ozx
1GAOll+J8saUyB5qB4Vvh2Y8tMDeGJPGCd0bfq9nH7zebkiPvTCF1/lH6Yzj47K4
mLIHKcWfZfNHIgE/T8YtnWFYi4O6mAq7m8UH6jtBnnpfh79TqBe5rZtDLPzebmcz
X0p1bZbAqNcmCDMEw+VOf2w7JV/zYz8Fat9z50K+DDy1v9e/eScBtRHs1BNJR2LO
mqPKTgrQruDn6SzHtQcL3+IQ6uazJixv8869zyhRgYu7lh+ZArD00tH3KYLmAdnB
eo/vM3k6qbiv56mB0TtUuIN2TGThegyYFiOa+AS4AVpDp3XcSzo/YeO9g/urCPvx
0PdWJIr1PZjsSNuCnO/R7kdoDwhNVnxtY4rcXBgX4bIW0dHlUgjgVIzDNQeSrBIO
UvcstvXZ+2YGLQwkilXN1zzLMevY5F4K6+K3btkjBO735lJA7pXtodlsrZtUu/de
SLD0KLphbx1RMOVtXZ96KH9hmGlYCADAygI7Ip59TIGI2p6O6oUK7wxO72RA+poO
e4nIDC4E/oFHoJhOgHsOwD/EUPXgW1gKXt3mx8Tj9cdkfiaWb5Jf16dhoZvDQF2I
EKFkWSd+Ey9afUwEoiwTfvWS91O2i6l/m+KMjIKEOgnuxpN+2YM9mgdlD79DHWOt
DRZJgxmSjzgrCdQtdZukQtR8r7ye6az9csf39N1h4v8oD/nOPj30+HyiHX/7AT7I
Z0XmLZ00j69S528NGy3J7QWHXStfOFl2wHrLceO0viamxMD7eg7ZUgmrYDXGtC/Z
QYUCK/LmW1mRMXO8al60ahRfIYzS2epaKNxNsZyjiWk4zOQOxBgOog+l47Ok/dK4
1oMGX9EfmKo3w4NHsLux2PZebv40DImOYH0253fFULkDYH+04EEx4C17irnUDiJK
Y7inx+Bc0wJTTeg0Oa6DPogqjB1SnDOahERT7ZMGrBZscHEaDBsYmM/1N5pPcjK1
/WDOWpxiny6o4Z+jlDh4YXOyJeqtAN2Z659GysLuPsqRSHM3FcjtqbvOCyyrkIIi
x9djIym+6LlBA7WnA/aArfXR/Lr/wljXfneKy21ulyQ8xylc3g+xnjQq/29QpqNY
hqHngLS+4ykTiMdoV0C8ikI6S2V3J9HA37fysqEYq3v+urRMP2bgHurjgemiKpX9
E0zYtFOtrp0bS75kCOMl/ELQVFnKTkmWreA7Btjagy6r3ro0LJgc7L4WNzq4RefZ
7AmdlnY2rSIcqyUIApKWy6XjleAgVTr+wrYYy5xCsl3rRabLMNGFbS3XQ6fwgKDA
bXOqL7iGxClkdMde7WpoZMfXuO10V/S/yhpbq3hDi8sbEp5VvAVkRnuV585ZHW94
+nxGLOIP3L1X8+C+6BvcTSr8+HdCsfb01JSnZmTQA0ac6HU4MGJW4ApfUocm4/Db
GI5Hl2DFQV1AguViLcscs5LHEO3GBw+KiiJxYa1Zm4MQ8DfwWLDuqjxnTYcLRckY
PIgFEGC0oZDdltW5tCGMz6ViCBsv94Ev4RWLx3mNFGOMnRNiql1f+p5UZ3qHDMLn
ErojdlSEkrDZaLiCgJRH3aa4NvY7hWVhvexgH4ogQLv+1ANXD7qfceTvI3HDlbbz
Zqb2T9C7aElQ/BvQ2S49ajcJmw+lH4LEn7TDw5Hsz2Q2htWvOZ7m/TxiTWOTDoNw
ChuJKdBDEKpT8WvTkcjoQeftr1bmHiS37zCFN22IlbTmikub8u7c2/0OPzhqO1CQ
r15unVEE2R6synnpX2gvrknG++en6d5ExlxwGCFjvJ4QHIDDXRe5twgTJkhdmZmK
NVQ1RHITlu6BLRTCXImlG1JsSi3PQEmfofQEMlPSpkIgLr6/ApGyFxXO/LdA9iGa
mYEWzzicvJOAlwNA314HE+mk/7548BGu/a6tNFkYYlQ16ZgWfE+Ow/JlyVoCBsqy
mANnh2vOu+KW5N9Bm7q/RNWIgES/G8XQbwXvP1dFxQFG4DCGmjCYW52409HxEWfb
r0nvD10ZiHf4ej70g6JXmkcDT9Zp48uf2V6snxhoUEfPPO117QujtrJo5p08sgCV
dKsGJHWzDJLHsHan5jOUlkG8ZxqO1MRyJ/lks1xy32a0BcTcAgH4h6sOzc1c5Hgc
8967Kbmf8+IY6xC4J38XSpbmlg/oVtpUqG8PLMMSC5SphQhOE4qqplIuIJD3YOkS
uPKaYcnZYSrC0nbo+WW73n3stqCJBqZ5TPRSY8TSw5gwB9PskiQ1KiciQJox+gHm
GhDyjilnc88b+axGn8epvxkgWc0WUoB+q/cCqOiEpqZImJDFfKeoACYVqI14/fPG
3h1B065Z7+sbA0EiRhQmYnxSjtE+m4ahU2BcIk2tgFCg3JwPFKkGA8LqQaez9/tb
nOFLcS0Hf/FmdLq6WzKeNmiEfVKBlEcPFpeN8vEGz1KKG5jZtfE6qOhHkQ4smdFD
kxFJPmlxnT+GvTr4UxNKPr32SuaSzX7T8Z+VPKeZoR2rOC16pZNUxxucpWtCvpDQ
lv6F32cT1NyvzYC0yYKKADVzt1HJE5MVa71GOZw8o2YEk6EAan5xpF1SXMW/XgsH
R8hwKxr/AvTq1qN3B5BtUDpIfX1qJX9gDflIxElZW/KaEOaRV5SfHSVa1lzl2At6
ZWmwuv9nBUvbZWlAAnx202CG7low3LmZgtFAmU32S4ydPcNAEmWa43D5KUyOZgHm
7yjP7K4jsFyzc5cm5Wcq+2+w5uq0A3eKyFRWMKnYcaY9u4sMELR9lflCpf/x8KeG
oI461r9rs83pRNRFuKc8mZNYJYSd5+WfYeTKPK435jkONwj2HdDH7GmTvCOITTmJ
xexYkQe3NuhzP/uCCd43u/dR0Ynk9ZwC80qTfDoGJBAPuhxOW0/tREvlv+QEVeZt
1zCM9GRXdJ4HaxY9uUuo9PAMVvgC3HEVujC63xgqDl8fH2s+A+yK7eZDrsESdRtv
92qqf8RGMRJDqPazIbC+3Q6oneS8OEYZSn2c2z2xVD1qcmzasX/blwIaxihY985/
ISWNUowDCSgykSwU8RzfnfCOMWfiKmbUxGU+hzCN8GADBoGctPAoTfv3aRAhGmdw
u4SiRf8uzG18P6hghly35ghJgcP1uqfeekduFq8vdS015akczbVBzoTn0/wMFyrK
aQk1fo4ISTStpAF6QmRVqdfjJNtSRJ7fAV03uuid3xHjVzRc+ZIiwtJJaJT1WivO
164sEHx3IenVmVnK2fD4IbDpZG8PCyeqrcjnIpMfNSAyedkot88ktmqGX6nDhKTz
HOFkj13GksF6Yroo7gwd1XujYsT1lPxdzobtnA45sb9gn7AqbUFrPZpWspgChifW
dNQ9fc7LZlPbNd0CXqKpj/RYz4TPm7LDHN8uePP+JgIZFWX2zLPRn26RRpuQWoes
FVBJFXP3+kigG3s8GpYgYSTRdq1mFnzrMnxgk1mJqWT6NJ6BPw8FgGB+3A6PfzfS
X8qthvq3x8cDklmk0paECgcExKqahIaNce7gK7VwlZjmmAZ6U8wCPAaWGOF/KqvX
CXJhCpl0UB3GtNkOkDF2yWOBjPyao++9kM6ZyYjGsrDA7a/tLmAZ36j4ZboUzX3x
Di4WnzQvKH5ACeB/j/G5062/o35ZX8h1JgZZjskQ8mhl0ZKF8dPVBtPWmjyws0/v
G2dNC47aOCi9MmR16VqNqF5hQpT3Kc76gQXcyyfYf+cLCeVOb9WdNx6CD9f26hsy
hegSBXV/fMj99acNF59sGM2wczqZVDSzSbqGknV6dN9j3HQFIClDpENtMni/UbHB
UUxLDTEUqK54BlEECf5JAW2PVBfbk4QfmX5xpkvW/AUz1+eZaZfp5FYZ45bp3LBU
ibFXLLaTjlbSpEGGsVU0/2qeKyDLnxxWW17x56gO7T6ALHbHyyyyCEc4bvumu3a3
ekhMpDHDYG4rWVu/OARHRZ4TeZL35xMlpB0lVBwVWhc8LnjDq4NPc8Rqr5b3yrl8
eb5Qo6ictvHK1o95cKWNSKDTJggvJj+iG0nKQJTc9snJR04aChbH4MSOAhCeDtX1
fOjVqko1YtHD2ZL68kKo4cqQgx99DDCgKdlEdHuDtj2y4p33+yb0qm7ZcgwhD41C
JWzaXtwMXgOfj++6cEKdu59ZKWelBdkgb/XSYrojiwRRmyOhceg1J4upEJaBDFcw
c0dbPqyTKYbddgamN34XQ05LcJaP/TxtRknvxuuh7OPsy0x6ZHQMEDUvGzymr1eM
99jEedbE39vzH/ktzYrwQq+rPn3dVvp8Fwy3wFHRtOpZBBsPaIiEUnn87TAzqP6w
TZNqffWSR2vQk2GW0YhCEkrgxVyL4RUCZF8q0nrxUR9AwXndic/2Nserwz0IMZ54
MujEoZGlUwMgcIfucDT9SFVDVHlrWxHZ1fEByKX+WKIuXzM2TH4x8+x7oc3787pU
cm15bmSg7f+LgpJWsGpsOM+PwYq2W2T3oYAR+yhNs2t7EZ1/RUbeych7F+sAcOY+
86nRO/e05PgD/d/u7S3HoSmjWC7qw2ioYatJOmGWI+kY+ZgqI3p50utx8OsjXj0L
0X/gwsyucxoE4YW8sSxrR7e6XyfaqE1ORlO/N2xuAuI0sptHtGPwKfZwd3IcruiF
/1oLwP1FcMzXkuMR4GfLjP/LUHdNlY8OmIA3qVChzYJgh3BRF+m6xUu3AGQjfZnu
MPlsz55dwfV3AY/YIT644nIhQfm4GWt93HSNI5/QJA2tIDWFLcoiFxNkHOz+yvvK
wOK+GPCESExqrmdh/McMCJxNX2RReUUSYPOwIl8HPQ5K4EIa4yVgKgue1i/wxvim
vZ06DTOI4jQLRuW4gj6wk7xKDg+iN0wLIsMb2Sf+uqdV0q2QPySPnfWYOiMBTcyx
SeTvxgDWFmPIon8DEh+RVFCQqQ5rtUzCxWb5mjpaQnhbeljC/ZKn1VedRBXFoVL4
umPBKnwJ9jlgE5wAH/lKEwow9GO68fmOcnJYt0G2sECSSSytr0KhmQS0BXs2jrMu
Zuax3rzQrDzfa3WbuCsjLac2GR0k5DxxEYDe3DB3KTKbqnw/4anUHB7SRx6Pbp8A
znmgi+o9IeffCOAD6EmmgcW6rh8dz65us6ENAXHiig9LT0PbgzxZVmsRVcJQhSGJ
2pfGLZ9t23Ohu6u/y6pi6fmAV1MnPpszE4HMHmBs5j7XjHK4FBak3jga05f46RPV
MSavphxLJaWMKp+WEOuwEj8gQq8D2LDrySOq57A6d2Nq9ctRVXsas1xW788ck4hZ
NU+6tyK5rnHn8gXowqwi4GFq+RHyKmmATG3iGplqrAiFpINrMNP6z1eMo4C7iGBg
W+tfv7pqzp5IxVIH1UMIUuv7GMlw0Wt/6805x+XIC9iiHIz52xD28/dPb9IDsUAd
hshTezWrFHV6B1o6FDI47mtbMDEbv88ahz1IbHL4EYVa4JElaKEDxHX81Pt6KdwP
0oowWhRIBPhcivEOvvqdTLtV2CsCWmVMGu1SX+mSCNBUDl1F0GkboeW5ckZoftAs
b5RgewRftIeMS2B3oMpcKF1eGE1xvas8bqo6SsG8DmLqNXuylW/SaRfk8n1C2X1e
+WEIIXHcwGnjIhHC+EOEVewrpd+xriLBIDi4aeqrnxHBUlLdn6vLlwnzJDCaVGw8
+fuLOyWFil9hVJVzViftrrIWhykWQ2yTI0EEHG/dPVe/eKEIlfOoLalqkCUl2YUO
W+PZIEQ1SlNsupPeG9u3FcdDCBPNzjEMw9sGMoiWROcvepNYTep1l75zxAJvVRqX
eULDVLZuDciT6+m6X5mQoorlMATp/f6o69o+mK8OE1AYjc/MGIG4aGPQI8sMmnXN
3cpp2+p2yKTiWHdH+5clfFWlzQmE9OImLtP+A2Rn74Z920Aujv694UQtLA+gikLc
fs2DUuXZAkyUp4yRg5RhzVXeWnYwmBjq0D3Vqpfkn0ZcfOcOr7qXHYjLztf+msZA
d8hkgSiJ5nOiJvC3sbw72oMO5LiQwEVLdacFOkw9WCAqoSWc+boUMJrUyHXaN9V1
B6Rd8xfqF7mcZ796VPdxLWsXSkSrERmy+sQY+ZF+qvqPl2RRjT9dy8qIPJtVxWig
IilJEOm0tKaWFO9Jcn/xW5B7+NQUlvzxZbE/SzCf1/BSpwoogXNPyXXX3t+HpzsW
UroWk6EqB1rEdO4fdLjBr8Mk6G1eXbrnHWxVmmPuT+2aiY/wTjqubN4fUvst2aTp
jiUQpXaysqneJJrBxgRJ+GFju3Nquw2RC3SAQBMjX0pd2WpTXZnttkHv7A8mgozj
dtQghQS1qLaLedg5XBpDiOXzLSzXwuzfVN2iMzsj6vN9JWIP42how4RNiUsHOLpS
yUTd1TXsT0dgt28aZO+P69KAXU7Jguv8Yq48l6gzujg43T8nVpCI/ML4y/EpnrfB
yOZ5zX6cpqbLdcH5lhw4j01uRioV7HcidJF46BGOpfnGKUcFt9Nry1vrrO3VDSvb
n3GNnUyTWb5D6DSKeD4wRT38FQ7sD28nzANoF/OUFq9bXLFbOlqaLHHUZT/mD4Xy
mInbgxRNIc6QYwOmgwCLfS2SldFXWFO4ikp0pg2FCIL4w2m9i+JbQKeT5I3OuEfr
30q2rLRDd+aRfb3FQD76ffwyL8MjzfXsiXq1LcAMCs5DD5mkZ4io3HClF+fMScfB
HEF6ctpp1S6FL/yDDfWdAUw9v1ooliVWuN0MemO1/5QWZFOcobAKZtCQgTL0fXfd
vcSn0t2bNyEsrYgEeglhVH5awKDYODX7iHmrIkwmkLYPAgFJrYx6IOflWcHxE0Xj
wM0IQVEXrmdtQ6KuTDa6Qr5dWLqdGTcWuZ2ezzjuOz3WznwNHir2GQK6VFPd410e
EzD/baS9onnbwc3X0wAxnsW/nIAXcLU0i4u5XFuQY86inEjA8XS0IGIKavEJRIjk
Upuj20JYug/UEX/UxEsJdVz1VUTumKPZyqJD5jxeT5Oi0IyvSM4KcUIrrGA2vhjJ
/Tz8o2tGIoeAtXREW9GHua1KGtVvD52da7Q5Q8Kpd5JCgwp8sP7cB2hgPKHeA2CU
ETJgxX4eWikZvTPfzscaT33DDtTz2Ngn73ZPtmN8uwqN9I59kfQEK4qJB+n5H6BZ
DoJgR/TytgvRtCG0BLf1tYSnXOcY8dB/M3iaKF7O8oMAZAiTiFeuZgW8VytTav9U
l+qvYkVQbcM8tLEN6LDIozU/Aa/54eohtovPOOBjCxj4/QVBTTr7i5QpeheyF466
BwVEZOObJJGQjBSu925NkvARmjL6LY3lQujEpBl92r0B5p57K6ZfXdIM6+2phokQ
toPr5BCuhNZgjxl26tk6cwJYxmJHqzvJmCUYcIOtkUWqDQDK09tOtno9IuW+THOX
RElKZ8QtZVpl+lQ0RREEVy1XHrEI0LWKPWBPOEV+ZQThA3IG+RZFRI8asNPcnRx6
1yU4xXoJ38KHidsyROnVGvJX88BgE1edN1ORqDTilLzhYdwdvSUiSaUBqBXCknjw
3GRGSPqnqfH5Og7uIPjiFfvIHtG53mhJD51uqmEAmHvsOrXRLF4bFdAWYikc4GaZ
uWjE9v6CLfrxVSJAH24n1Wq40YJRl0WUlR6vhjayu5UyluCuGfzHt7kgMUfeQ7ei
R7eRn0LPSt4ivE0XG6KYtQiDQfXyuDc4tfs8ug9W6x7F91Rqldtz1eHg1NYIfoHQ
yXuLvuNba3tNJViEOj8feN2kvyq6BR/6JwzSMUc4mm6uimK/RLldIRjMMRBTYAZl
qulerL5LsqeP22zXMK7LG/iFkcB+PKzf249M83tWJbXIvP0ZqK2//xyEtbh5LGfW
FT72zcYVNwp4Bsu+/7W0eRg0epBLk535OlX6UCkNsNuSXeoD1f3QbswQhqL47eWk
e4x4ZbH9vRqVbBQdHw3uN8Qj2k7oKNx9FtwT5Ogi/QxIpuU7PdNjwpD8qkiQ641Z
Ban2R3oinTMU3SCTkhqc9QMcw5r0N1AUtI4T+xaE5EyQXIXxZ41dItR9mS0EYgcU
7335qsQbvayM8myT9iiLnjGtbD5tWph2d2cL2Wyah58IWWjwA00xSVFPoLg+VM3l
9uKoDpMLsJU42DfMQCPF5FMKhTYESpWtnTEsyaKyXxvuicEsvdkNFM8GXlMqHmZ7
yhv5qTsoo8HJxHzCCuPIS6AozghMp0+sSuT5+HijjhX7Tum1zHBly/J5S7R+IBq0
HuH2Lw3gyz0zz7jUIw2Ou83nT45cwiIP20ELDduayE4fRjcAJQaiUvVIr5fv7bVM
vYhe3zHc0n/4EAzxh4oScTe4siB6OzENu6DxkZK9Vrmd8whUA+3bHTcGmMH9exPd
utbQX+l9YC0q4JFuGD8M5G6VLQgtDhAQuGS/yPs42YXYzStJWp5sdCp2lA2XkekP
fRFGEFEBB65RYWKtNsXRzUPpGFn5Pj4INvsmaz+5ywYBcJqWG7dlQwFIXXW+pP+P
iJp88E3fOtLclfMsH6ReSQ/qSfjP/9AGhY6nXSlhuaL1ynbH0dEF4+asR3FgrHhd
z/Ju+8Lw41yNVnC404QBxXds4XGzcgDRdhE8cR0h9cg6zLIDSC/FZKymSzK9mGh0
lUjuDxPmkz20ZzN4u5ddr88JqMxhpY4JFu6GLXzb+PVDp15X26qliek4gSz24j3f
2rqDeYy8zpMP/jVSrEx4oi4AhMIVWQWLVMp9Hah3PqvgaVaSoavqe8CtWUsmtHNn
Wm0fNkQpV0ppKtzUxsltMzMd1MAlUutfH/J6r0JFne7E0spNiHlLeC2KBAaqWKoQ
Xmh+YgfVUv+IuLzZWBDzwIBw7k/TYXGLLlCzZhSOF5wAwX8zTMMfDhgs3hTxJkwY
i2z8ZZgjEbrOlSgblBI2HeDNLRrdlNMVhD7xHVU2L3Ojuez9KLaCoBsKgbR9t2ZX
sY+tGJul9V5ZSqwhLnsB3kakIcxv261wh+YGgZElNj8Ug89gNliQ0cGHalI7lttK
OXrH5safwYmTAQOiIhdtlX/pUnrqKTbTF1Fhk17TACwsVSjnCpEPe3Vx4EpKOtLu
sHK7IbOC2lJ32bWtFeDhqSpxHiPM81MV2nW2hyoatg5SQ2bXLlbLm51J/1KoOLhX
NT4bUnoHf/t4kAaN7VaPupSbq39GtOcxHvYiwxNNzwpVLDEx+ib09/Xzdq2g2hoW
DXbyR4CsmIzP191kD6t19nk9mcaPfeJ4uJXAK1Q+BNvrLy+pO8oc0I+kKI/TDxjR
Df8ejfeY/MS+BCCujWTpWjwfeIaAkLPsqUG+yImzJuK02CrirNek/i0LAAto2G2V
xL4ySWfmPXqDJrH1MxaY7VkFcLORZ8NPbok9eyAC28Ek4ZaPM4HA28V5GxvELEvg
fizHGwsBB3teouaZgyh2hRKOsJ+Td1Smt8cLjYiMTC0lmWyxZstPW7KFdTTrfsXR
z5m3bNaqDEtVaE1neGorYTid8505qfmgEK83fH1acR48/WlfUVQDXFifXzAXtOHK
x8ily6Mu4gchR9/BMGntk85bYdH6ZJUS4W4AzU40DR8vXQ0btwC3x6nX/93iMtAZ
i8sqlcKd88lAGRDSq14HcQpzThtl0MdoLn/t+Nfm7ZNCGM/2bc5XZiBczyZ/gF+Y
CYTAgYGvuS0UqM24xrLTDl0JwE1DIstWhiUAUEyx3MrQD3YxgsYI6K93dJ/gLRPo
d4yL3H588clkbSrCxn8ZMdQK2oyLj3r0Ccf/J2BGT4P2NEheXW0wZk2z6oywl5Xl
zPKCA65eoa9J9go8KUpiZyPRIUNGHHalKWw9jWscg/PBRZ+LDa+ZA9yVU9UUDc3k
ofO8d+19Ouey7hJ+/y5UIyZKnLMZBgyr3nZ7pyK3vjGg78j+QGmfd/8RNTnj8g6+
87HHu7p6yH5Wyzt/1VZNkoMmCrfolcBtr5NGIz1Cp+PJZg+wKYL+lGaxNvl1WQeB
a9QUkZjHi7wDPshdlZiWR4crs/XNmj4em2l7G1bEVPCV6m7ZsorljqirCqX9L2Eg
hcoee0GUB8YluId8N9d/0LQnCqnVC4g2Bsu08Xtjl4+KkhWiT3gRLoA5vJLyV14K
hfeI0BkzU8VKR7AycGvOICzL17sAKN0EJvaqlNXfY5ouV41Q/sfSUNu0yLIyuPwN
4gWqbcDiRa2RPUVME9HJ161p7Uz/whgAXKzN5v9gSBFSOqYAa61ArDe9j/9CUrRf
WXf+WGHDP/ieBIHNOksFGPGIal7ENP28vKYaBNKEJWnNTciDyeXYp2nsD5KTlm2D
CyBsbr5V4YSAyWszcSH0uwgMYxQ00CVEgHz7QJj3mQb7lsNOcDTk/N4S2AFdIzhB
ayX2LbmMfIJPYMNBU4pcorlqEItE7S0UNe/gIcapLeOalsUrPopuY/Y8jKRFr6eK
iOLV/4cLp31U4GTOmyrbr61QgTJeZkeP7YgW2WAEruXmUhA0Fwqpbd8TZ3gQzZEw
+SGS/BCoQJBz3C1iiMHHnRMmCm7Z8tRAXSvUYlHtgB9+hv/BJaJayPvaesmQGsIS
T8r98HeIPTVGR+yaSdnBE2Qykh0ki74JugNTOlROk2YfSyCnroni9hCMRWHxOH1P
yHbnjNLlpgZP6J3Cpy1vaf7SXASDMRM1yvCF5urpIIln7Dyr/ttkMK9RRzPhFLYB
A5o40BFYyToqa8+v7hjfN38YFYuXDmmZt16+dBHrEgsQiPrAXVh8jWBs3TrlVhlE
UHmNrkKC9HtLeQzLk/WpQEOeWAcSBaah74wDLZjV2Agpe7tJ30sGvvww5yGGIY5M
CNeHiNRiVhRXcs+1NiSQ4/dHUvM8koR4opesRRmSnotreSbA61O3IxaKyM0wu16B
q2wP7Vx0NldfWOKfQYCzT71xFTpb62wZs7tz6yx29k21xmBaunxsWgyHaVZc7V2s
PHpIDuXDtM7DzARAH6Vi7kCdlTbDbmBFmbEYNrFIQYKj1OkGLfBqaVARn1He5Aj/
BpEpJRk8h9EpjJo9taHYW9o8tcOUnfWHZ0uHW/BqszcyjtzC9Gw+Yw4V8+ucbnwE
ximlF3QYoexXtXL8pBo3MwO8ebiV8Ky+mvtQe0pVDn2hg0wI1OEAHKw0gEs4NA9L
ptY8VaC34XEC6Bt29coUyTOzy2fpueIWkRYrnGQTTh5firpzq0LStu0NfZsk38Pl
/j6vnqXLdYiPLrqV+cWcUcoTMDbffg7BQinPabO2gIm/0j+GWtUvvqQbH3Y+5gan
rwQcAWJrptH/r8ZRuhp4U3IINpWAfUH3SDYAkWKdtMQY5VGmvLaBpV6Sjy3VMgkO
QDzImYbGQ5NtonexlY+GZpB+/DAdQ9bWSqCxxLzwW1bIK5+1q0dmCItEvYZY/+LI
reBaoWO09sQEatpb35br5Zy34Vz1+xUb9a8YTWATwpB56keXcmmWPn0oF6dTE0Pq
iPcPPDnvfh8nFY5XmBJXVGhNUzLkB59NppU5s9rZSvb757w1vj8qxTbAQI8EHifE
ipnAH5B3pJ69ZwHsRfxRVMTbpGf5m3AKSnfl0tUsu2kpZ8ZOFLPoxW3Yy45B3TQQ
MfUgf2SvJ9ugs4LZv96GdlVz0K8c7hG2MjGlN4DWDEK+8nL4SCBbr4UzbK3tMpx/
vkrRSz7aE4DIqQ4Bw2It40wRL+lCSTgDiNijl1SOQkwxb+dgVxhSfs8iDx+19/3C
8ilNWSmTLs2KHOdzh4XpI0HUxyhAdudvAxVomaNVAKzpTg1C8i8cWol0YSNeeyvN
9un7BfvXKJtUngJqExY+90WF3rq4K5H8Y/XJkQoGeVLDx1lo4BlisKZyeagmPCPq
musKWgyRBj3gYpNiS1MBDr+osbeWD6wR0Ynlre8Fno25TpC4IfmqXuexZKngF2Dr
zixS+xq4Pvj4ubFfs4kC/4zausOuNlFZWx1ShsM/Zlsd5QClJVb1yOIwBd0fyHIW
RUFhIe1CQNzxXdjemmRw7Vyx4VxVHfjQiZBtzN0cOrwWQ5WbOtV91Zz8JVCiHF+s
SD96ajh7T4fvKX2FADcbOvS+44abIfILbmv/8kqh1CAksT9E3z10Y4mGSk76U0vn
lpYMe2dpBDaKTgq3LIiIlEjpPh8u1JnN9IS1v7DteYe08I+t7qjtO/htbJJtQtT0
BD6qm8dkfqiYNhD6omiRaYZmUfcq/zN12VDmoSy28dodALA1v6BQUP2Nr1sO3y2s
qdBSyOwzXAgFCaQeP7cVt4fXappVkuqdS4GswSrgxYD0D0L902glJbCFofEvhUPg
7heJRwFt96Tt1GEh8l0F3F4y9p9HkIrQjV6v1G895sOd4rY37jCTi0UT+wjcLtWQ
OtB3zDXG6ljjkAJ3EwK/SFKFIkag2QHKj1e4Bh0A23mvKpYSgmWKch2jh++tFwPp
RBLTp3kYVciy24q/ema7+hZZoo3ki58u9PyNYmxA0slmGY7FHyzY8hh1exNbSCnC
+or7YOgfNoQ4bk0bxlcOko27TKe+efyRyMpwMKmuW5W8ntFcwa8k+x+JLvwqAyMa
7tpnjcm6JLY7lA+vCCT3QqGQ8kNMjZopd5bT6GkeLlpQAm2v4IgQh2tmJh9rkW+F
STGRVzPuUH01uhgho/hHbNfAgaG3Hy/9QkHs+6tfbTEXmM+5CZI38ulb5o0OWgMR
c8rxpd8b17JYIpbPwsee2Uud4eKVGgeLPaLQRrbMMLr28uf5MEjOcy1Inq/O1gey
OixU9B30JFWEqSuJf96cpSxvzE+IAjD+aLAv3+K/yQCtkElfyPpshN469i2RjQAf
w7j9FqbDWgRNpwP+aj3vxDIRjgUEHyBO7uxJHertUyozqzkHAfLkaWc1UZTrOFxA
8fKQ559OVuVENbxNY23Nm806tL60am4d7UPNOB3036Y8ZuE63XQAwUtl/vnT72+M
O5XBl6W1wImE7V2fREczJx0os0Dm8R0oLnFToC9A6Fs419jIMS7e63efEb0TLC0R
625dLM50aTeHkWFnqvqwr6UDfWhqQ5Wg+8tvL9S38rszFHIdOlV8kvcik38L/1d4
PF2CQbo1K0aONIrA5Inha8UKfssE8Y3KBurdVirQuzm1y/ibFqd/JyxJBepmI0ok
iqsLd0Pd5TX66q7p/V7UHYCh4mF08A+Oo7yaU77GyLg0Yr0MHwxzBzhfH07B03vG
L96Zh6lES5lhA60MMyvp0gEIZZHJCNXM0e1pEb5DhC0K4FwykeW76q/LDGpoL//z
Vw/RhMF9oLOO/TFh8UhaIoIkjl3Kyr9IAKfvgdVUvC4wTMulx/mNLM0/uLMJTDWz
K+ZFuw1cMu4JF5tNGoAcELYF6dPsTdmzHyMQZP16WyApiEkzkZpBv6Bsq958Q2rj
hiqrdpoXUfkPunIlEqMKf4a0fjp7qNXL/x8zyUgupF7FzPVD3zSZKWuBuFKU7Oqj
uPFsqECT5oVvQIv1j0mO+ce+zw8vgL9QKn4VnauEvO/qYEinGi2Lr38NTgklU0hR
hDRq3F3+ihLcJ6W2vPWH1lR6ChZDQuoj+kfomHEgJn0PzzwDtSyTbfZODw6Nt2nL
H94fr8SPuyQOs8Moi60vpXOZpjZz4GO/JfqY+0MLA7T8fR5AFWVyQfoZzQXfTx4e
aHzJ3R0ngQgz+HX2HIlnU4MRQ7f9Oacsn1DH0CygUdZ3QU0k5JlqZxv4do8HqK4P
RAYxQWHqPsmpGKNWeauZlieHqIKyv1+p071Fox3GcfqTJoHNsfazS6+5fAlerxMo
Ka3WSO9lBa25nCPG7gGLdbP3UpTGl6e3o709R7IPGbEoqfPp0Nm9woyoOfHDQrl5
lGbB1KjP8DJ+R7qNx6Yu282f9KUTpi+QkEYjY17jFHaKQV3jOZnA6m4ybcY5dh8k
Ls5VnkbA3iTxVbRBuLMwfsiy8g6Unk4Mkld337Ha+pieMifXs/yOLlB6bc2+j+w1
0eikPxjo3mawK+2xtEgwGpmFjOvqaSeIGN3VDLKgn+RflM31VwUmq4k9nMYuXmjw
oAUATLh26VDGN3gkCbwzGSgyvIgdlsBEiSuVmrf23DwECUFnPGhXF/3uKh327EZC
wxYcrI6em98PdIM2IzKovV1NqR5t+BeDJQczd6VLdHmDFl6VeLuLCyYeSsbtkkwr
t/2Wqh1PYd8N9CY/X1boTR/D5qsQTbCKumvFD15JafqWVmeEEHJI3mfPrSzNdQqt
3OCLQaw+TkOAM+R/H+/t39yZShM9yyyQNqlCFQg7R8ZoWBX8fJTqRjFZGZoUsm/f
fOsBH4sJ83upoxCOU1oFCKxNt/Wt3pq65z2Y5LIrx4TN0Ln6Z62IemrvE/hIYdfv
hqpTwLM08MvP+E46Z65/T7Rvw+Rm1vafJ0gvPOgGnxhE+OFI7d2Qh95nBwkzXyiu
qKd4gAVn4pmv118aUSuTSaH9tcUoGtA0jezYlQztgWCR1VzddfoYGjzFrHSDH1hL
eJjGqVJTx6POijX7ckj7AiKFvGWcWosr38NwytySJTXEiY1GTtgYu3JolbZxwa7e
9ZBnvSLGAX9ILngLgmVcxxhPFnl30mB0gPBKFQcc6R08wlPrnKroygUypl0YxnxQ
5AC0hGD+Es6KDPcfwToSrMdwfONsh8vdui6MQMgS33IqtjlPkDZ6hPMM85i6Iuwp
m9A7E88oSvjc6/q51AbIbYAc0i+IV4MSN27ssTwHfI1ub4NbaYHDeYtbvEIUC7Sv
zL2E0FwkdMFld/47UI49S2yngoa1MOspc8rnkvbBxdUSlcj4wBj7BSZYtK/83Av7
ujkWdujfS8Eu27KbCyWpgrIRCaPdB9UGz1goeyVtEIziJ0efMIdoQ+W2o57SpkbU
vEXBGuXGUTTzLGR5ne0+ZFbzpgw9iluj5SHrEbvCs/xpkn1r1Eg5u9pvelqRKu65
IYWEqOjlBf7shiYOmgM7wrLjkw9a2W9LL+n3xXmsgct9WnQ1hFeLl22IT/53K/Lm
2pGEnfZXs3JLDSNGrBEb0t6VKtfgfzChpUSzpRAi8bWSJm08a5C1VaXCjZAsN4i4
XrS6BMSAiXQdo1ReuOPjraHE569QF5msAtEvFpfhZoNUEWuRB6LSJ4oJkIFtuNJy
N5J2iMU2LtqsB3vMxh+SIG+paidu55I6GF6+KZA0kXVxnPHf/XMQFdeIF2ezorJj
TGBQx8cTtbTuHdXEphw6pftxw65nA2dd1gbXG4FeYkFnfZtNGwy7RitbSXrHsFvY
EiH8VSoaRhiExrvnPFNRTlE/pUOEkx68mAk8bmYEv9+dSW5D5/j0hWGNzN71iAGL
LWXTIEAFmEUMvbxCcTbovu1r5BMKPeeO70EcPg/ZSFvheP7fjQ+/1Tik0FBBKjLV
e/K8erP0rg65CaZMuUqNFGlay65yur99dOsE8PklN0aeYdXuZyF2h8ByRWddO+f/
`pragma protect end_protected
